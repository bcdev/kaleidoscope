netcdf PE_mro_mean_error_prv_4km_120p_spring_cor {
dimensions:
	lat = 4320 ;
	lon = 8640 ;
variables:
	float latitude(lat) ;
		latitude:_FillValue = -999.f ;
		latitude:units = "degrees north" ;
		latitude:_Storage = "contiguous" ;
		latitude:_Endianness = "little" ;
	float longitude(lon) ;
		longitude:_FillValue = -999.f ;
		longitude:units = "degrees east" ;
		longitude:_Storage = "contiguous" ;
		longitude:_Endianness = "little" ;
	double alphaB(lat, lon) ;
		alphaB:_FillValue = -999. ;
		alphaB:units = "mgC mgChl-1 h-1 (W m-2)-1" ;
		alphaB:_Storage = "contiguous" ;
		alphaB:_Endianness = "little" ;
	double PmB(lat, lon) ;
		PmB:_FillValue = -999. ;
		PmB:units = "mgC mgChl-1 h-1" ;
		PmB:_Storage = "contiguous" ;
		PmB:_Endianness = "little" ;
	double lat(lat) ;
		lat:_FillValue = NaN ;
		lat:_Storage = "contiguous" ;
		lat:_Endianness = "little" ;
	double lon(lon) ;
		lon:_FillValue = NaN ;
		lon:_Storage = "contiguous" ;
		lon:_Endianness = "little" ;
	double alphaB_unc(lat, lon) ;
		alphaB_unc:_FillValue = -999. ;
		alphaB_unc:units = "mgC mgChl-1 h-1 (W m-2)-1" ;
		alphaB_unc:_Storage = "contiguous" ;
		alphaB_unc:_Endianness = "little" ;
	double PmB_unc(lat, lon) ;
		PmB_unc:_FillValue = -999. ;
		PmB_unc:units = "mgC mgChl-1 h-1" ;
		PmB_unc:_Storage = "contiguous" ;
		PmB_unc:_Endianness = "little" ;

// global attributes:
		:description = "Physio_parameters_spring" ;
		:source = "netCDF3 python" ;
		:history = "Created Thu Jul  4 09:47:53 2024" ;
		:_NCProperties = "version=2,netcdf=4.9.2,hdf5=1.14.3" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
}
