netcdf \200001-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0-1M {
dimensions:
	lat = 3600 ;
	lon = 7200 ;
	time = 1 ;
variables:
	float lat(lat) ;
		lat:_FillValue = NaNf ;
		lat:standard_name = "latitude" ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
		lat:actual_range = -89.975f, 89.975f ;
		lat:axis = "Y" ;
		lat:reference_datum = "geographical coordinates, WGS84 projection" ;
		lat:comment = "Latitude geographical coordinates, WGS84 projection" ;
		lat:bounds = "lat_bnds" ;
		lat:_Storage = "chunked" ;
		lat:_ChunkSizes = 3600 ;
		lat:_Shuffle = "true" ;
		lat:_DeflateLevel = 1 ;
		lat:_Endianness = "little" ;
	float lon(lon) ;
		lon:_FillValue = NaNf ;
		lon:standard_name = "longitude" ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
		lon:actual_range = -179.975f, 179.975f ;
		lon:axis = "X" ;
		lon:reference_datum = "geographical coordinates, WGS84 projection" ;
		lon:comment = "Longitude geographical coordinates, WGS84 projection" ;
		lon:bounds = "lon_bnds" ;
		lon:_Storage = "chunked" ;
		lon:_ChunkSizes = 7200 ;
		lon:_Shuffle = "true" ;
		lon:_DeflateLevel = 1 ;
		lon:_Endianness = "little" ;
	float analysed_sst(time, lat, lon) ;
		analysed_sst:_FillValue = NaNf ;
		analysed_sst:long_name = "analysed sea surface temperature" ;
		analysed_sst:standard_name = "sea_water_temperature" ;
		analysed_sst:units = "kelvin" ;
		analysed_sst:valid_min = -300s ;
		analysed_sst:valid_max = 4500s ;
		analysed_sst:actual_range = 271.15f, 305.09f ;
		analysed_sst:source = "ATSR<1,2>-ESACCI-L3U-v3.0, AATSR-ESACCI-L3U-v3.0, SLSTR<A,B>-ESACCI-L3U-ICDR-v3.0 AVHRR<06,07,08,09,10,11,12,14,15,16,17,18,19>_G-ESACCI-L3U-v3.0, AVHRRMT<A,B>-ESACCI-L3U-v3.0, AMSR<E,2>-ESACCI-L2P-v2.0" ;
		analysed_sst:depth = "20 cm" ;
		analysed_sst:ancillary_variables = "analysed_sst_uncertainty mask" ;
		analysed_sst:_Storage = "chunked" ;
		analysed_sst:_ChunkSizes = 1, 1800, 3600 ;
		analysed_sst:_Shuffle = "true" ;
		analysed_sst:_DeflateLevel = 4 ;
		analysed_sst:_Endianness = "little" ;
	float analysed_sst_uncertainty(time, lat, lon) ;
		analysed_sst_uncertainty:_FillValue = NaNf ;
		analysed_sst_uncertainty:long_name = "estimated error standard deviation of analysed_sst" ;
		analysed_sst_uncertainty:standard_name = "sea_water_temperature standard_error" ;
		analysed_sst_uncertainty:units = "kelvin" ;
		analysed_sst_uncertainty:valid_min = 0s ;
		analysed_sst_uncertainty:valid_max = 32767s ;
		analysed_sst_uncertainty:actual_range = 0.11f, 2.86f ;
		analysed_sst_uncertainty:ancillary_variables = "mask" ;
		analysed_sst_uncertainty:_Storage = "chunked" ;
		analysed_sst_uncertainty:_ChunkSizes = 1, 1800, 3600 ;
		analysed_sst_uncertainty:_Shuffle = "true" ;
		analysed_sst_uncertainty:_DeflateLevel = 4 ;
		analysed_sst_uncertainty:_Endianness = "little" ;
	float sea_ice_fraction(time, lat, lon) ;
		sea_ice_fraction:_FillValue = NaNf ;
		sea_ice_fraction:long_name = "sea ice area fraction" ;
		sea_ice_fraction:standard_name = "sea_ice_area_fraction" ;
		sea_ice_fraction:units = "1" ;
		sea_ice_fraction:valid_min = 0b ;
		sea_ice_fraction:valid_max = 100b ;
		sea_ice_fraction:actual_range = 0.f, 1.f ;
		sea_ice_fraction:source = "EUMETSAT_OSI-SAF-ICE-OSI-450, EUMETSAT_OSI-SAF-ICE-OSI-430-b" ;
		sea_ice_fraction:comment = " Sea ice area fraction" ;
		sea_ice_fraction:ancillary_variables = "mask" ;
		sea_ice_fraction:_Storage = "chunked" ;
		sea_ice_fraction:_ChunkSizes = 1, 1800, 3600 ;
		sea_ice_fraction:_Shuffle = "true" ;
		sea_ice_fraction:_DeflateLevel = 4 ;
		sea_ice_fraction:_Endianness = "little" ;
	float mask(time, lat, lon) ;
		mask:_FillValue = NaNf ;
		mask:standard_name = "status_flag" ;
		mask:long_name = "sea/land/lake/ice field composite mask" ;
		mask:valid_min = 1b ;
		mask:valid_max = 31b ;
		mask:actual_range = 1b, 14b ;
		mask:flag_masks = 1b, 2b, 4b, 8b, 16b ;
		mask:flag_meanings = "water land optional_lake_surface sea_ice optional_river_surface" ;
		mask:source = "Carrea, L.; Embury, O.; Merchant, C.J. (2015): GloboLakes: high-resolution global limnology dataset v1. Centre for Environmental Data Analysis, 21 July 2015. doi:10.5285/6be871bc-9572-4345-bb9a-2c42d9d85ceb (described in: Carrea, L., Embury, O. and Merchant, C. J. (2015) Datasets related to in-land water for limnology and remote sensing applications: distance-to-land, distance-to-water, water-body identifier and lake-centre co-ordinates. Geoscience Data Journal, 2 (2). pp. 83-97. doi:10.1002/gdj3.32), Schaffer, J.; Timmermann, R. (2016): Greenland and Antarctic ice sheet topography, cavity geometry, and global bathymetry (RTopo-2), links to NetCDF files. PANGAEA, doi:10.1594/PANGAEA.856844 (supplement to: Schaffer, J.; Timmermann, R.; Arndt, J.E.; Kristensen, S.S.; Mayer, C.; Morlighem, M.; Steinhage, D. (2016): A global, high-resolution data set of ice sheet topography, cavity geometry, and ocean bathymetry. Earth System Science Data, 8(2), 543-557, doi:10.5194/essd-8-543-2016)" ;
		mask:comment = "b0: 1=grid cell is open sea water b1: 1=grid cell is land b2: 1=grid cell is lake surface b3: 1=grid cell is sea ice b4-b7: reserved for future grid mask data" ;
		mask:_Storage = "chunked" ;
		mask:_ChunkSizes = 1, 1800, 3600 ;
		mask:_Shuffle = "true" ;
		mask:_DeflateLevel = 4 ;
		mask:_Endianness = "little" ;
	int time(time) ;
		time:long_name = "reference time of sst field" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:comment = "" ;
		time:bounds = "time_bnds" ;
		time:units = "seconds since 1970-01-01" ;
		time:calendar = "proleptic_gregorian" ;
		time:_Storage = "contiguous" ;
		time:_Endianness = "little" ;

// global attributes:
		:Conventions = "CF-1.5, Unidata Observation Dataset v1.0" ;
		:title = "ESA SST CCI Analysis v3.0" ;
		:summary = "European Space Agency Sea Surface Temperature Climate Change Initiative: Analysis product version 3.0" ;
		:references = "Embury, O. et al. Satellite-based time-series of sea-surface temperature since 1980 for climate applications. Scientific Data (2024). https://doi.org/10.1038/s41597-024-03147-w" ;
		:institution = "ESACCI" ;
		:history = "Created using OSTIA reanalysis system CDR3.0. Composite generated by NEODAAS using weighted mean equal to sum(analysed_sst / (analysed_sst_uncertainty**2)) / sum(1/(analysed_sst_uncertainty**2)). Composite using: 20000101120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000102120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000103120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000104120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000105120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000106120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000107120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000108120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000109120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000110120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000111120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000112120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000113120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000114120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000115120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000116120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000117120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000118120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000119120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000120120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000121120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000122120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000123120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000124120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000125120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000126120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000127120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000128120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000129120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000130120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc, 20000131120000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-GLOB_CDR3.0-v02.0-fv01.0.nc" ;
		:comment = "These data were produced at the Met Office as part of the ESA SST CCI project. WARNING Some applications are unable to properly handle signed byte values. If values are encountered > 127, please subtract 256 from this reported value. Subsetting and compositing by NEODAAS" ;
		:license = "Creative Commons Attribution 4.0 https://creativecommons.org/licenses/by/4.0/ \n",
			"Users of these data should cite the dataset along with the dataset paper: Embury, O. et al. Satellite-based time-series of sea-surface temperature since 1980 for climate applications. Scientific Data (2024). https://doi.org/10.1038/s41597-024-03147-w" ;
		:id = "OSTIA-ESACCI-L4-GLOB_CDR-v3.0" ;
		:naming_authority = "org.ghrsst" ;
		:product_version = "3.0.1" ;
		:uuid = "92fbdb08-855d-4eb1-bb74-ae8c7a184405" ;
		:tracking_id = "92fbdb08-855d-4eb1-bb74-ae8c7a184405" ;
		:gds_version_id = "2.0" ;
		:netcdf_version_id = "4.3.2" ;
		:date_created = "20211125T002143Z" ;
		:file_quality_level = 3 ;
		:spatial_resolution = "0.05 degree" ;
		:start_time = "20000101T000000Z" ;
		:time_coverage_start = "20000101T000000Z" ;
		:stop_time = "20000201T000000Z" ;
		:time_coverage_end = "20000201T000000Z" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_resolution = "P1D" ;
		:source = "ATSR<1,2>-ESACCI-L3U-v3.0, AATSR-ESACCI-L3U-v3.0, SLSTR<A,B>-ESACCI-L3U-ICDR-v3.0 AVHRR<06,07,08,09,10,11,12,14,15,16,17,18,19>_G-ESACCI-L3U-v3.0, AVHRRMT<A,B>-ESACCI-L3U-v3.0, AMSR<E,2>-ESACCI-L2P-v2.0, EUMETSAT_OSI-SAF-ICE-OSI-450-v2.0, EUMETSAT_OSI-SAF-ICE-OSI-430-b" ;
		:platform = "ERS-<1,2>, Envisat, Sentinel-3<A,B>, NOAA-<06,07,08,09,10,11,12,14,15,16,17,18,19>, MetOp<A,B>, Aqua, GCOM-W" ;
		:sensor = "ATSR, AATSR, SLSTR, AVHRR, AMSR" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:metadata_link = "https://doi.org/10.5285/4a9654136a7148e39b7feb56f8bb02d2" ;
		:doi = "10.5285/4a9654136a7148e39b7feb56f8bb02d2" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = 0.05f ;
		:geospatial_lon_min = -180.f ;
		:geospatial_lon_max = 180.f ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = 0.05f ;
		:northernmost_latitude = 90.f ;
		:southernmost_latitude = -90.f ;
		:easternmost_longitude = 180.f ;
		:westernmost_longitude = -180.f ;
		:geospatial_vertical_min = -0.2f ;
		:geospatial_vertical_max = -0.2f ;
		:acknowledgment = "The European Space Agency (ESA) funded the research and development of software to generate these data (grant reference ESA/AO/1-9322/18/I-NB), in addition to funding the production of the Climate Data Record (CDR) for 1980 to 2021. The Copernicus Climate Change Service (C3S) funded the development of the Interim-CDR (ICDR) extension and production of ICDR during 2022. From 2023 onwards the production of the ICDR is funded by the UK Natural Environment Research Council (NERC grant reference number NE/X019071/1, Earth Observation Climate Information Service) and the UK Marine and Climate Advisory Service (UKMCAS), benefitting from the Earth Observation Investment Package of the Department of Science, Innovation and Technology." ;
		:creator_name = "Met Office" ;
		:creator_url = "https://www.metoffice.gov.uk" ;
		:creator_email = "ml-ostia@metoffice.gov.uk" ;
		:creator_type = "institution" ;
		:creator_institution = "Met Office" ;
		:project = "Climate Change Initiative - European Space Agency" ;
		:contributor_name = "JASMIN" ;
		:contributor_role = "This work used JASMIN, the UK\'s collaborative data analysis environment (https://jasmin.ac.uk)" ;
		:publisher_name = "NERC EDS Centre for Environmental Data Analysis" ;
		:publisher_url = "https://www.ceda.ac.uk" ;
		:publisher_email = "support@ceda.ac.uk" ;
		:publisher_type = "institution" ;
		:processing_level = "L4" ;
		:cdm_data_type = "grid" ;
		:product_specification_version = "SST_CCI-PSD-UKMO-201-Issue-2" ;
		:key_variables = "analysed_sst,sea_ice_fraction" ;
		:contact = "https://climate.esa.int/en/projects/sea-surface-temperature" ;
		:citation = "If you use this data towards any publication, please acknowledge NEODAAS in addition to ESA using: \'The authors thank the NERC Earth Observation Data Acquisition and Analysis Service (NEODAAS) for supplying data for this study\' and then email NEODAAS (info@neodaas.ac.uk) with the details. The service relies on users\' publications as one measure of success." ;
		:_NCProperties = "version=2,netcdf=4.8.1,hdf5=1.12.1" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 0 ;
		:_Format = "netCDF-4 classic model" ;
}
