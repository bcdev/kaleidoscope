netcdf ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1M_MONTHLY_4km_GEO_PML_OCx_QAA-200001-fv6.0 {
dimensions:
	time = 1 ; // was UNLIMITED (1 currently)
	lat = 4320 ;
	lon = 8640 ;
variables:
	float Rrs_412(time, lat, lon) ;
		Rrs_412:_FillValue = 9.96921e+36f ;
		Rrs_412:ancillary_variables = "Rrs_412_rmsd Rrs_412_bias" ;
		Rrs_412:long_name = "Sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 412 nm." ;
		Rrs_412:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFV13N26" ;
		Rrs_412:standard_name = "surface_ratio_of_upwelling_radiance_emerging_from_sea_water_to_downwelling_radiative_flux_in_air" ;
		Rrs_412:units = "sr-1" ;
		Rrs_412:units_nonstandard = "sr^-1" ;
		Rrs_412:wavelength = 412 ;
		Rrs_412:_Storage = "chunked" ;
		Rrs_412:_ChunkSizes = 1, 270, 270 ;
		Rrs_412:_Shuffle = "true" ;
		Rrs_412:_DeflateLevel = 3 ;
		Rrs_412:_Endianness = "little" ;
	float Rrs_412_bias(time, lat, lon) ;
		Rrs_412_bias:long_name = "Bias of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 412 nm." ;
		Rrs_412_bias:_FillValue = 9.96921e+36f ;
		Rrs_412_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_bias.dat" ;
		Rrs_412_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_412_bias:rel = "uncertainty" ;
		Rrs_412_bias:units = "sr-1" ;
		Rrs_412_bias:units_nonstandard = "sr^-1" ;
		Rrs_412_bias:wavelength = 412 ;
		Rrs_412_bias:_Storage = "chunked" ;
		Rrs_412_bias:_ChunkSizes = 1, 270, 270 ;
		Rrs_412_bias:_Shuffle = "true" ;
		Rrs_412_bias:_DeflateLevel = 3 ;
		Rrs_412_bias:_Endianness = "little" ;
	float Rrs_412_rmsd(time, lat, lon) ;
		Rrs_412_rmsd:long_name = "Root-mean-square-difference of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 412 nm." ;
		Rrs_412_rmsd:_FillValue = 9.96921e+36f ;
		Rrs_412_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_rmsd.dat" ;
		Rrs_412_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_412_rmsd:rel = "uncertainty" ;
		Rrs_412_rmsd:units = "sr-1" ;
		Rrs_412_rmsd:units_nonstandard = "sr^-1" ;
		Rrs_412_rmsd:wavelength = 412 ;
		Rrs_412_rmsd:_Storage = "chunked" ;
		Rrs_412_rmsd:_ChunkSizes = 1, 270, 270 ;
		Rrs_412_rmsd:_Shuffle = "true" ;
		Rrs_412_rmsd:_DeflateLevel = 3 ;
		Rrs_412_rmsd:_Endianness = "little" ;
	float Rrs_443(time, lat, lon) ;
		Rrs_443:_FillValue = 9.96921e+36f ;
		Rrs_443:ancillary_variables = "Rrs_443_rmsd Rrs_443_bias" ;
		Rrs_443:long_name = "Sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 443 nm." ;
		Rrs_443:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFV13N26" ;
		Rrs_443:standard_name = "surface_ratio_of_upwelling_radiance_emerging_from_sea_water_to_downwelling_radiative_flux_in_air" ;
		Rrs_443:units = "sr-1" ;
		Rrs_443:units_nonstandard = "sr^-1" ;
		Rrs_443:wavelength = 443 ;
		Rrs_443:_Storage = "chunked" ;
		Rrs_443:_ChunkSizes = 1, 270, 270 ;
		Rrs_443:_Shuffle = "true" ;
		Rrs_443:_DeflateLevel = 3 ;
		Rrs_443:_Endianness = "little" ;
	float Rrs_443_bias(time, lat, lon) ;
		Rrs_443_bias:long_name = "Bias of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 443 nm." ;
		Rrs_443_bias:_FillValue = 9.96921e+36f ;
		Rrs_443_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_bias.dat" ;
		Rrs_443_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_443_bias:rel = "uncertainty" ;
		Rrs_443_bias:units = "sr-1" ;
		Rrs_443_bias:units_nonstandard = "sr^-1" ;
		Rrs_443_bias:wavelength = 443 ;
		Rrs_443_bias:_Storage = "chunked" ;
		Rrs_443_bias:_ChunkSizes = 1, 270, 270 ;
		Rrs_443_bias:_Shuffle = "true" ;
		Rrs_443_bias:_DeflateLevel = 3 ;
		Rrs_443_bias:_Endianness = "little" ;
	float Rrs_443_rmsd(time, lat, lon) ;
		Rrs_443_rmsd:long_name = "Root-mean-square-difference of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 443 nm." ;
		Rrs_443_rmsd:_FillValue = 9.96921e+36f ;
		Rrs_443_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_rmsd.dat" ;
		Rrs_443_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_443_rmsd:rel = "uncertainty" ;
		Rrs_443_rmsd:units = "sr-1" ;
		Rrs_443_rmsd:units_nonstandard = "sr^-1" ;
		Rrs_443_rmsd:wavelength = 443 ;
		Rrs_443_rmsd:_Storage = "chunked" ;
		Rrs_443_rmsd:_ChunkSizes = 1, 270, 270 ;
		Rrs_443_rmsd:_Shuffle = "true" ;
		Rrs_443_rmsd:_DeflateLevel = 3 ;
		Rrs_443_rmsd:_Endianness = "little" ;
	float Rrs_490(time, lat, lon) ;
		Rrs_490:_FillValue = 9.96921e+36f ;
		Rrs_490:ancillary_variables = "Rrs_490_rmsd Rrs_490_bias" ;
		Rrs_490:long_name = "Sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 490 nm." ;
		Rrs_490:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFV13N26" ;
		Rrs_490:standard_name = "surface_ratio_of_upwelling_radiance_emerging_from_sea_water_to_downwelling_radiative_flux_in_air" ;
		Rrs_490:units = "sr-1" ;
		Rrs_490:units_nonstandard = "sr^-1" ;
		Rrs_490:wavelength = 490 ;
		Rrs_490:_Storage = "chunked" ;
		Rrs_490:_ChunkSizes = 1, 270, 270 ;
		Rrs_490:_Shuffle = "true" ;
		Rrs_490:_DeflateLevel = 3 ;
		Rrs_490:_Endianness = "little" ;
	float Rrs_490_bias(time, lat, lon) ;
		Rrs_490_bias:long_name = "Bias of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 490 nm." ;
		Rrs_490_bias:_FillValue = 9.96921e+36f ;
		Rrs_490_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_bias.dat" ;
		Rrs_490_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_490_bias:rel = "uncertainty" ;
		Rrs_490_bias:units = "sr-1" ;
		Rrs_490_bias:units_nonstandard = "sr^-1" ;
		Rrs_490_bias:wavelength = 490 ;
		Rrs_490_bias:_Storage = "chunked" ;
		Rrs_490_bias:_ChunkSizes = 1, 270, 270 ;
		Rrs_490_bias:_Shuffle = "true" ;
		Rrs_490_bias:_DeflateLevel = 3 ;
		Rrs_490_bias:_Endianness = "little" ;
	float Rrs_490_rmsd(time, lat, lon) ;
		Rrs_490_rmsd:long_name = "Root-mean-square-difference of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 490 nm." ;
		Rrs_490_rmsd:_FillValue = 9.96921e+36f ;
		Rrs_490_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_rmsd.dat" ;
		Rrs_490_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_490_rmsd:rel = "uncertainty" ;
		Rrs_490_rmsd:units = "sr-1" ;
		Rrs_490_rmsd:units_nonstandard = "sr^-1" ;
		Rrs_490_rmsd:wavelength = 490 ;
		Rrs_490_rmsd:_Storage = "chunked" ;
		Rrs_490_rmsd:_ChunkSizes = 1, 270, 270 ;
		Rrs_490_rmsd:_Shuffle = "true" ;
		Rrs_490_rmsd:_DeflateLevel = 3 ;
		Rrs_490_rmsd:_Endianness = "little" ;
	float Rrs_510(time, lat, lon) ;
		Rrs_510:_FillValue = 9.96921e+36f ;
		Rrs_510:ancillary_variables = "Rrs_510_rmsd Rrs_510_bias" ;
		Rrs_510:long_name = "Sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 510 nm." ;
		Rrs_510:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFV13N26" ;
		Rrs_510:standard_name = "surface_ratio_of_upwelling_radiance_emerging_from_sea_water_to_downwelling_radiative_flux_in_air" ;
		Rrs_510:units = "sr-1" ;
		Rrs_510:units_nonstandard = "sr^-1" ;
		Rrs_510:wavelength = 510 ;
		Rrs_510:_Storage = "chunked" ;
		Rrs_510:_ChunkSizes = 1, 270, 270 ;
		Rrs_510:_Shuffle = "true" ;
		Rrs_510:_DeflateLevel = 3 ;
		Rrs_510:_Endianness = "little" ;
	float Rrs_510_bias(time, lat, lon) ;
		Rrs_510_bias:long_name = "Bias of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 510 nm." ;
		Rrs_510_bias:_FillValue = 9.96921e+36f ;
		Rrs_510_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_bias.dat" ;
		Rrs_510_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_510_bias:rel = "uncertainty" ;
		Rrs_510_bias:units = "sr-1" ;
		Rrs_510_bias:units_nonstandard = "sr^-1" ;
		Rrs_510_bias:wavelength = 510 ;
		Rrs_510_bias:_Storage = "chunked" ;
		Rrs_510_bias:_ChunkSizes = 1, 270, 270 ;
		Rrs_510_bias:_Shuffle = "true" ;
		Rrs_510_bias:_DeflateLevel = 3 ;
		Rrs_510_bias:_Endianness = "little" ;
	float Rrs_510_rmsd(time, lat, lon) ;
		Rrs_510_rmsd:long_name = "Root-mean-square-difference of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 510 nm." ;
		Rrs_510_rmsd:_FillValue = 9.96921e+36f ;
		Rrs_510_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_rmsd.dat" ;
		Rrs_510_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_510_rmsd:rel = "uncertainty" ;
		Rrs_510_rmsd:units = "sr-1" ;
		Rrs_510_rmsd:units_nonstandard = "sr^-1" ;
		Rrs_510_rmsd:wavelength = 510 ;
		Rrs_510_rmsd:_Storage = "chunked" ;
		Rrs_510_rmsd:_ChunkSizes = 1, 270, 270 ;
		Rrs_510_rmsd:_Shuffle = "true" ;
		Rrs_510_rmsd:_DeflateLevel = 3 ;
		Rrs_510_rmsd:_Endianness = "little" ;
	float Rrs_560(time, lat, lon) ;
		Rrs_560:_FillValue = 9.96921e+36f ;
		Rrs_560:ancillary_variables = "Rrs_560_rmsd Rrs_560_bias" ;
		Rrs_560:long_name = "Sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 560 nm." ;
		Rrs_560:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFV13N26" ;
		Rrs_560:standard_name = "surface_ratio_of_upwelling_radiance_emerging_from_sea_water_to_downwelling_radiative_flux_in_air" ;
		Rrs_560:units = "sr-1" ;
		Rrs_560:units_nonstandard = "sr^-1" ;
		Rrs_560:wavelength = 560 ;
		Rrs_560:_Storage = "chunked" ;
		Rrs_560:_ChunkSizes = 1, 270, 270 ;
		Rrs_560:_Shuffle = "true" ;
		Rrs_560:_DeflateLevel = 3 ;
		Rrs_560:_Endianness = "little" ;
	float Rrs_560_bias(time, lat, lon) ;
		Rrs_560_bias:long_name = "Bias of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 560 nm." ;
		Rrs_560_bias:_FillValue = 9.96921e+36f ;
		Rrs_560_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_bias.dat" ;
		Rrs_560_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_560_bias:rel = "uncertainty" ;
		Rrs_560_bias:units = "sr-1" ;
		Rrs_560_bias:units_nonstandard = "sr^-1" ;
		Rrs_560_bias:wavelength = 560 ;
		Rrs_560_bias:_Storage = "chunked" ;
		Rrs_560_bias:_ChunkSizes = 1, 270, 270 ;
		Rrs_560_bias:_Shuffle = "true" ;
		Rrs_560_bias:_DeflateLevel = 3 ;
		Rrs_560_bias:_Endianness = "little" ;
	float Rrs_560_rmsd(time, lat, lon) ;
		Rrs_560_rmsd:long_name = "Root-mean-square-difference of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 560 nm." ;
		Rrs_560_rmsd:_FillValue = 9.96921e+36f ;
		Rrs_560_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_rmsd.dat" ;
		Rrs_560_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_560_rmsd:rel = "uncertainty" ;
		Rrs_560_rmsd:units = "sr-1" ;
		Rrs_560_rmsd:units_nonstandard = "sr^-1" ;
		Rrs_560_rmsd:wavelength = 560 ;
		Rrs_560_rmsd:_Storage = "chunked" ;
		Rrs_560_rmsd:_ChunkSizes = 1, 270, 270 ;
		Rrs_560_rmsd:_Shuffle = "true" ;
		Rrs_560_rmsd:_DeflateLevel = 3 ;
		Rrs_560_rmsd:_Endianness = "little" ;
	float Rrs_665(time, lat, lon) ;
		Rrs_665:_FillValue = 9.96921e+36f ;
		Rrs_665:ancillary_variables = "Rrs_665_rmsd Rrs_665_bias" ;
		Rrs_665:long_name = "Sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 665 nm." ;
		Rrs_665:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFV13N26" ;
		Rrs_665:standard_name = "surface_ratio_of_upwelling_radiance_emerging_from_sea_water_to_downwelling_radiative_flux_in_air" ;
		Rrs_665:units = "sr-1" ;
		Rrs_665:units_nonstandard = "sr^-1" ;
		Rrs_665:wavelength = 665 ;
		Rrs_665:_Storage = "chunked" ;
		Rrs_665:_ChunkSizes = 1, 270, 270 ;
		Rrs_665:_Shuffle = "true" ;
		Rrs_665:_DeflateLevel = 3 ;
		Rrs_665:_Endianness = "little" ;
	float Rrs_665_bias(time, lat, lon) ;
		Rrs_665_bias:long_name = "Bias of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 665 nm." ;
		Rrs_665_bias:_FillValue = 9.96921e+36f ;
		Rrs_665_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_bias.dat" ;
		Rrs_665_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_665_bias:rel = "uncertainty" ;
		Rrs_665_bias:units = "sr-1" ;
		Rrs_665_bias:units_nonstandard = "sr^-1" ;
		Rrs_665_bias:wavelength = 665 ;
		Rrs_665_bias:_Storage = "chunked" ;
		Rrs_665_bias:_ChunkSizes = 1, 270, 270 ;
		Rrs_665_bias:_Shuffle = "true" ;
		Rrs_665_bias:_DeflateLevel = 3 ;
		Rrs_665_bias:_Endianness = "little" ;
	float Rrs_665_rmsd(time, lat, lon) ;
		Rrs_665_rmsd:long_name = "Root-mean-square-difference of sea surface reflectance defined as the ratio of water-leaving radiance to surface irradiance at 665 nm." ;
		Rrs_665_rmsd:_FillValue = 9.96921e+36f ;
		Rrs_665_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/rrs/cci_Rrs_rmsd.dat" ;
		Rrs_665_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		Rrs_665_rmsd:rel = "uncertainty" ;
		Rrs_665_rmsd:units = "sr-1" ;
		Rrs_665_rmsd:units_nonstandard = "sr^-1" ;
		Rrs_665_rmsd:wavelength = 665 ;
		Rrs_665_rmsd:_Storage = "chunked" ;
		Rrs_665_rmsd:_ChunkSizes = 1, 270, 270 ;
		Rrs_665_rmsd:_Shuffle = "true" ;
		Rrs_665_rmsd:_DeflateLevel = 3 ;
		Rrs_665_rmsd:_Endianness = "little" ;
	float adg_412(time, lat, lon) ;
		adg_412:_FillValue = 9.96921e+36f ;
		adg_412:ancillary_variables = "adg_412_rmsd adg_412_bias" ;
		adg_412:long_name = "Absorption coefficient for dissolved and detrital material at 412 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		adg_412:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		adg_412:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		adg_412:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		adg_412:units = "m-1" ;
		adg_412:units_nonstandard = "m^-1" ;
		adg_412:wavelength = 412 ;
		adg_412:_Storage = "chunked" ;
		adg_412:_ChunkSizes = 1, 270, 270 ;
		adg_412:_Shuffle = "true" ;
		adg_412:_DeflateLevel = 3 ;
		adg_412:_Endianness = "little" ;
	float adg_412_bias(time, lat, lon) ;
		adg_412_bias:long_name = "Bias of absorption coefficient for dissolved and detrital material at 412 nm." ;
		adg_412_bias:_FillValue = 9.96921e+36f ;
		adg_412_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_bias.dat" ;
		adg_412_bias:ref = "http://www.uncertweb.org" ;
		adg_412_bias:rel = "uncertainty" ;
		adg_412_bias:units = "m-1" ;
		adg_412_bias:units_nonstandard = "m^-1" ;
		adg_412_bias:wavelength = 412 ;
		adg_412_bias:_Storage = "chunked" ;
		adg_412_bias:_ChunkSizes = 1, 270, 270 ;
		adg_412_bias:_Shuffle = "true" ;
		adg_412_bias:_DeflateLevel = 3 ;
		adg_412_bias:_Endianness = "little" ;
	float adg_412_rmsd(time, lat, lon) ;
		adg_412_rmsd:long_name = "Root-mean-square-difference of absorption coefficient for dissolved and detrital material at 412 nm." ;
		adg_412_rmsd:_FillValue = 9.96921e+36f ;
		adg_412_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_rmsd.dat" ;
		adg_412_rmsd:ref = "http://www.uncertweb.org" ;
		adg_412_rmsd:rel = "uncertainty" ;
		adg_412_rmsd:units = "m-1" ;
		adg_412_rmsd:units_nonstandard = "m^-1" ;
		adg_412_rmsd:wavelength = 412 ;
		adg_412_rmsd:_Storage = "chunked" ;
		adg_412_rmsd:_ChunkSizes = 1, 270, 270 ;
		adg_412_rmsd:_Shuffle = "true" ;
		adg_412_rmsd:_DeflateLevel = 3 ;
		adg_412_rmsd:_Endianness = "little" ;
	float adg_443(time, lat, lon) ;
		adg_443:_FillValue = 9.96921e+36f ;
		adg_443:ancillary_variables = "adg_443_rmsd adg_443_bias" ;
		adg_443:long_name = "Absorption coefficient for dissolved and detrital material at 443 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		adg_443:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		adg_443:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		adg_443:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		adg_443:units = "m-1" ;
		adg_443:units_nonstandard = "m^-1" ;
		adg_443:wavelength = 443 ;
		adg_443:_Storage = "chunked" ;
		adg_443:_ChunkSizes = 1, 270, 270 ;
		adg_443:_Shuffle = "true" ;
		adg_443:_DeflateLevel = 3 ;
		adg_443:_Endianness = "little" ;
	float adg_443_bias(time, lat, lon) ;
		adg_443_bias:long_name = "Bias of absorption coefficient for dissolved and detrital material at 443 nm." ;
		adg_443_bias:_FillValue = 9.96921e+36f ;
		adg_443_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_bias.dat" ;
		adg_443_bias:ref = "http://www.uncertweb.org" ;
		adg_443_bias:rel = "uncertainty" ;
		adg_443_bias:units = "m-1" ;
		adg_443_bias:units_nonstandard = "m^-1" ;
		adg_443_bias:wavelength = 443 ;
		adg_443_bias:_Storage = "chunked" ;
		adg_443_bias:_ChunkSizes = 1, 270, 270 ;
		adg_443_bias:_Shuffle = "true" ;
		adg_443_bias:_DeflateLevel = 3 ;
		adg_443_bias:_Endianness = "little" ;
	float adg_443_rmsd(time, lat, lon) ;
		adg_443_rmsd:long_name = "Root-mean-square-difference of absorption coefficient for dissolved and detrital material at 443 nm." ;
		adg_443_rmsd:_FillValue = 9.96921e+36f ;
		adg_443_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_rmsd.dat" ;
		adg_443_rmsd:ref = "http://www.uncertweb.org" ;
		adg_443_rmsd:rel = "uncertainty" ;
		adg_443_rmsd:units = "m-1" ;
		adg_443_rmsd:units_nonstandard = "m^-1" ;
		adg_443_rmsd:wavelength = 443 ;
		adg_443_rmsd:_Storage = "chunked" ;
		adg_443_rmsd:_ChunkSizes = 1, 270, 270 ;
		adg_443_rmsd:_Shuffle = "true" ;
		adg_443_rmsd:_DeflateLevel = 3 ;
		adg_443_rmsd:_Endianness = "little" ;
	float adg_490(time, lat, lon) ;
		adg_490:_FillValue = 9.96921e+36f ;
		adg_490:ancillary_variables = "adg_490_rmsd adg_490_bias" ;
		adg_490:long_name = "Absorption coefficient for dissolved and detrital material at 490 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		adg_490:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		adg_490:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		adg_490:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		adg_490:units = "m-1" ;
		adg_490:units_nonstandard = "m^-1" ;
		adg_490:wavelength = 490 ;
		adg_490:_Storage = "chunked" ;
		adg_490:_ChunkSizes = 1, 270, 270 ;
		adg_490:_Shuffle = "true" ;
		adg_490:_DeflateLevel = 3 ;
		adg_490:_Endianness = "little" ;
	float adg_490_bias(time, lat, lon) ;
		adg_490_bias:long_name = "Bias of absorption coefficient for dissolved and detrital material at 490 nm." ;
		adg_490_bias:_FillValue = 9.96921e+36f ;
		adg_490_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_bias.dat" ;
		adg_490_bias:ref = "http://www.uncertweb.org" ;
		adg_490_bias:rel = "uncertainty" ;
		adg_490_bias:units = "m-1" ;
		adg_490_bias:units_nonstandard = "m^-1" ;
		adg_490_bias:wavelength = 490 ;
		adg_490_bias:_Storage = "chunked" ;
		adg_490_bias:_ChunkSizes = 1, 270, 270 ;
		adg_490_bias:_Shuffle = "true" ;
		adg_490_bias:_DeflateLevel = 3 ;
		adg_490_bias:_Endianness = "little" ;
	float adg_490_rmsd(time, lat, lon) ;
		adg_490_rmsd:long_name = "Root-mean-square-difference of absorption coefficient for dissolved and detrital material at 490 nm." ;
		adg_490_rmsd:_FillValue = 9.96921e+36f ;
		adg_490_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_rmsd.dat" ;
		adg_490_rmsd:ref = "http://www.uncertweb.org" ;
		adg_490_rmsd:rel = "uncertainty" ;
		adg_490_rmsd:units = "m-1" ;
		adg_490_rmsd:units_nonstandard = "m^-1" ;
		adg_490_rmsd:wavelength = 490 ;
		adg_490_rmsd:_Storage = "chunked" ;
		adg_490_rmsd:_ChunkSizes = 1, 270, 270 ;
		adg_490_rmsd:_Shuffle = "true" ;
		adg_490_rmsd:_DeflateLevel = 3 ;
		adg_490_rmsd:_Endianness = "little" ;
	float adg_510(time, lat, lon) ;
		adg_510:_FillValue = 9.96921e+36f ;
		adg_510:ancillary_variables = "adg_510_rmsd adg_510_bias" ;
		adg_510:long_name = "Absorption coefficient for dissolved and detrital material at 510 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		adg_510:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		adg_510:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		adg_510:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		adg_510:units = "m-1" ;
		adg_510:units_nonstandard = "m^-1" ;
		adg_510:wavelength = 510 ;
		adg_510:_Storage = "chunked" ;
		adg_510:_ChunkSizes = 1, 270, 270 ;
		adg_510:_Shuffle = "true" ;
		adg_510:_DeflateLevel = 3 ;
		adg_510:_Endianness = "little" ;
	float adg_510_bias(time, lat, lon) ;
		adg_510_bias:long_name = "Bias of absorption coefficient for dissolved and detrital material at 510 nm." ;
		adg_510_bias:_FillValue = 9.96921e+36f ;
		adg_510_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_bias.dat" ;
		adg_510_bias:ref = "http://www.uncertweb.org" ;
		adg_510_bias:rel = "uncertainty" ;
		adg_510_bias:units = "m-1" ;
		adg_510_bias:units_nonstandard = "m^-1" ;
		adg_510_bias:wavelength = 510 ;
		adg_510_bias:_Storage = "chunked" ;
		adg_510_bias:_ChunkSizes = 1, 270, 270 ;
		adg_510_bias:_Shuffle = "true" ;
		adg_510_bias:_DeflateLevel = 3 ;
		adg_510_bias:_Endianness = "little" ;
	float adg_510_rmsd(time, lat, lon) ;
		adg_510_rmsd:long_name = "Root-mean-square-difference of absorption coefficient for dissolved and detrital material at 510 nm." ;
		adg_510_rmsd:_FillValue = 9.96921e+36f ;
		adg_510_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_rmsd.dat" ;
		adg_510_rmsd:ref = "http://www.uncertweb.org" ;
		adg_510_rmsd:rel = "uncertainty" ;
		adg_510_rmsd:units = "m-1" ;
		adg_510_rmsd:units_nonstandard = "m^-1" ;
		adg_510_rmsd:wavelength = 510 ;
		adg_510_rmsd:_Storage = "chunked" ;
		adg_510_rmsd:_ChunkSizes = 1, 270, 270 ;
		adg_510_rmsd:_Shuffle = "true" ;
		adg_510_rmsd:_DeflateLevel = 3 ;
		adg_510_rmsd:_Endianness = "little" ;
	float adg_560(time, lat, lon) ;
		adg_560:_FillValue = 9.96921e+36f ;
		adg_560:ancillary_variables = "adg_560_rmsd adg_560_bias" ;
		adg_560:long_name = "Absorption coefficient for dissolved and detrital material at 560 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		adg_560:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		adg_560:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		adg_560:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		adg_560:units = "m-1" ;
		adg_560:units_nonstandard = "m^-1" ;
		adg_560:wavelength = 560 ;
		adg_560:_Storage = "chunked" ;
		adg_560:_ChunkSizes = 1, 270, 270 ;
		adg_560:_Shuffle = "true" ;
		adg_560:_DeflateLevel = 3 ;
		adg_560:_Endianness = "little" ;
	float adg_560_bias(time, lat, lon) ;
		adg_560_bias:long_name = "Bias of absorption coefficient for dissolved and detrital material at 560 nm." ;
		adg_560_bias:_FillValue = 9.96921e+36f ;
		adg_560_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_bias.dat" ;
		adg_560_bias:ref = "http://www.uncertweb.org" ;
		adg_560_bias:rel = "uncertainty" ;
		adg_560_bias:units = "m-1" ;
		adg_560_bias:units_nonstandard = "m^-1" ;
		adg_560_bias:wavelength = 560 ;
		adg_560_bias:_Storage = "chunked" ;
		adg_560_bias:_ChunkSizes = 1, 270, 270 ;
		adg_560_bias:_Shuffle = "true" ;
		adg_560_bias:_DeflateLevel = 3 ;
		adg_560_bias:_Endianness = "little" ;
	float adg_560_rmsd(time, lat, lon) ;
		adg_560_rmsd:long_name = "Root-mean-square-difference of absorption coefficient for dissolved and detrital material at 560 nm." ;
		adg_560_rmsd:_FillValue = 9.96921e+36f ;
		adg_560_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_rmsd.dat" ;
		adg_560_rmsd:ref = "http://www.uncertweb.org" ;
		adg_560_rmsd:rel = "uncertainty" ;
		adg_560_rmsd:units = "m-1" ;
		adg_560_rmsd:units_nonstandard = "m^-1" ;
		adg_560_rmsd:wavelength = 560 ;
		adg_560_rmsd:_Storage = "chunked" ;
		adg_560_rmsd:_ChunkSizes = 1, 270, 270 ;
		adg_560_rmsd:_Shuffle = "true" ;
		adg_560_rmsd:_DeflateLevel = 3 ;
		adg_560_rmsd:_Endianness = "little" ;
	float adg_665(time, lat, lon) ;
		adg_665:_FillValue = 9.96921e+36f ;
		adg_665:ancillary_variables = "adg_665_rmsd adg_665_bias" ;
		adg_665:long_name = "Absorption coefficient for dissolved and detrital material at 665 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		adg_665:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		adg_665:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		adg_665:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		adg_665:units = "m-1" ;
		adg_665:units_nonstandard = "m^-1" ;
		adg_665:wavelength = 665 ;
		adg_665:_Storage = "chunked" ;
		adg_665:_ChunkSizes = 1, 270, 270 ;
		adg_665:_Shuffle = "true" ;
		adg_665:_DeflateLevel = 3 ;
		adg_665:_Endianness = "little" ;
	float adg_665_bias(time, lat, lon) ;
		adg_665_bias:long_name = "Bias of absorption coefficient for dissolved and detrital material at 665 nm." ;
		adg_665_bias:_FillValue = 9.96921e+36f ;
		adg_665_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_bias.dat" ;
		adg_665_bias:ref = "http://www.uncertweb.org" ;
		adg_665_bias:rel = "uncertainty" ;
		adg_665_bias:units = "m-1" ;
		adg_665_bias:units_nonstandard = "m^-1" ;
		adg_665_bias:wavelength = 665 ;
		adg_665_bias:_Storage = "chunked" ;
		adg_665_bias:_ChunkSizes = 1, 270, 270 ;
		adg_665_bias:_Shuffle = "true" ;
		adg_665_bias:_DeflateLevel = 3 ;
		adg_665_bias:_Endianness = "little" ;
	float adg_665_rmsd(time, lat, lon) ;
		adg_665_rmsd:long_name = "Root-mean-square-difference of absorption coefficient for dissolved and detrital material at 665 nm." ;
		adg_665_rmsd:_FillValue = 9.96921e+36f ;
		adg_665_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/adg/cci_iop_adg_rmsd.dat" ;
		adg_665_rmsd:ref = "http://www.uncertweb.org" ;
		adg_665_rmsd:rel = "uncertainty" ;
		adg_665_rmsd:units = "m-1" ;
		adg_665_rmsd:units_nonstandard = "m^-1" ;
		adg_665_rmsd:wavelength = 665 ;
		adg_665_rmsd:_Storage = "chunked" ;
		adg_665_rmsd:_ChunkSizes = 1, 270, 270 ;
		adg_665_rmsd:_Shuffle = "true" ;
		adg_665_rmsd:_DeflateLevel = 3 ;
		adg_665_rmsd:_Endianness = "little" ;
	float aph_412(time, lat, lon) ;
		aph_412:_FillValue = 9.96921e+36f ;
		aph_412:ancillary_variables = "aph_412_rmsd aph_412_bias" ;
		aph_412:grid_mapping = "crs" ;
		aph_412:long_name = "Phytoplankton absorption coefficient at 412 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		aph_412:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		aph_412:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		aph_412:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		aph_412:units = "m-1" ;
		aph_412:units_nonstandard = "m^-1" ;
		aph_412:wavelength = 412 ;
		aph_412:_Storage = "chunked" ;
		aph_412:_ChunkSizes = 1, 270, 270 ;
		aph_412:_Shuffle = "true" ;
		aph_412:_DeflateLevel = 3 ;
		aph_412:_Endianness = "little" ;
	float aph_412_bias(time, lat, lon) ;
		aph_412_bias:long_name = "Bias of phytoplankton absorption coefficient at 412 nm." ;
		aph_412_bias:_FillValue = 9.96921e+36f ;
		aph_412_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_bias.dat" ;
		aph_412_bias:ref = "http://www.uncertweb.org" ;
		aph_412_bias:rel = "uncertainty" ;
		aph_412_bias:units = "m-1" ;
		aph_412_bias:units_nonstandard = "m^-1" ;
		aph_412_bias:wavelength = 412 ;
		aph_412_bias:_Storage = "chunked" ;
		aph_412_bias:_ChunkSizes = 1, 270, 270 ;
		aph_412_bias:_Shuffle = "true" ;
		aph_412_bias:_DeflateLevel = 3 ;
		aph_412_bias:_Endianness = "little" ;
	float aph_412_rmsd(time, lat, lon) ;
		aph_412_rmsd:long_name = "Root-mean-square-difference of phytoplankton absorption coefficient at 412 nm." ;
		aph_412_rmsd:_FillValue = 9.96921e+36f ;
		aph_412_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_rmsd.dat" ;
		aph_412_rmsd:ref = "http://www.uncertweb.org" ;
		aph_412_rmsd:rel = "uncertainty" ;
		aph_412_rmsd:units = "m-1" ;
		aph_412_rmsd:units_nonstandard = "m^-1" ;
		aph_412_rmsd:wavelength = 412 ;
		aph_412_rmsd:_Storage = "chunked" ;
		aph_412_rmsd:_ChunkSizes = 1, 270, 270 ;
		aph_412_rmsd:_Shuffle = "true" ;
		aph_412_rmsd:_DeflateLevel = 3 ;
		aph_412_rmsd:_Endianness = "little" ;
	float aph_443(time, lat, lon) ;
		aph_443:_FillValue = 9.96921e+36f ;
		aph_443:ancillary_variables = "aph_443_rmsd aph_443_bias" ;
		aph_443:grid_mapping = "crs" ;
		aph_443:long_name = "Phytoplankton absorption coefficient at 443 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		aph_443:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		aph_443:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		aph_443:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		aph_443:units = "m-1" ;
		aph_443:units_nonstandard = "m^-1" ;
		aph_443:wavelength = 443 ;
		aph_443:_Storage = "chunked" ;
		aph_443:_ChunkSizes = 1, 270, 270 ;
		aph_443:_Shuffle = "true" ;
		aph_443:_DeflateLevel = 3 ;
		aph_443:_Endianness = "little" ;
	float aph_443_bias(time, lat, lon) ;
		aph_443_bias:long_name = "Bias of phytoplankton absorption coefficient at 443 nm." ;
		aph_443_bias:_FillValue = 9.96921e+36f ;
		aph_443_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_bias.dat" ;
		aph_443_bias:ref = "http://www.uncertweb.org" ;
		aph_443_bias:rel = "uncertainty" ;
		aph_443_bias:units = "m-1" ;
		aph_443_bias:units_nonstandard = "m^-1" ;
		aph_443_bias:wavelength = 443 ;
		aph_443_bias:_Storage = "chunked" ;
		aph_443_bias:_ChunkSizes = 1, 270, 270 ;
		aph_443_bias:_Shuffle = "true" ;
		aph_443_bias:_DeflateLevel = 3 ;
		aph_443_bias:_Endianness = "little" ;
	float aph_443_rmsd(time, lat, lon) ;
		aph_443_rmsd:long_name = "Root-mean-square-difference of phytoplankton absorption coefficient at 443 nm." ;
		aph_443_rmsd:_FillValue = 9.96921e+36f ;
		aph_443_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_rmsd.dat" ;
		aph_443_rmsd:ref = "http://www.uncertweb.org" ;
		aph_443_rmsd:rel = "uncertainty" ;
		aph_443_rmsd:units = "m-1" ;
		aph_443_rmsd:units_nonstandard = "m^-1" ;
		aph_443_rmsd:wavelength = 443 ;
		aph_443_rmsd:_Storage = "chunked" ;
		aph_443_rmsd:_ChunkSizes = 1, 270, 270 ;
		aph_443_rmsd:_Shuffle = "true" ;
		aph_443_rmsd:_DeflateLevel = 3 ;
		aph_443_rmsd:_Endianness = "little" ;
	float aph_490(time, lat, lon) ;
		aph_490:_FillValue = 9.96921e+36f ;
		aph_490:ancillary_variables = "aph_490_rmsd aph_490_bias" ;
		aph_490:grid_mapping = "crs" ;
		aph_490:long_name = "Phytoplankton absorption coefficient at 490 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		aph_490:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		aph_490:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		aph_490:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		aph_490:units = "m-1" ;
		aph_490:units_nonstandard = "m^-1" ;
		aph_490:wavelength = 490 ;
		aph_490:_Storage = "chunked" ;
		aph_490:_ChunkSizes = 1, 270, 270 ;
		aph_490:_Shuffle = "true" ;
		aph_490:_DeflateLevel = 3 ;
		aph_490:_Endianness = "little" ;
	float aph_490_bias(time, lat, lon) ;
		aph_490_bias:long_name = "Bias of phytoplankton absorption coefficient at 490 nm." ;
		aph_490_bias:_FillValue = 9.96921e+36f ;
		aph_490_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_bias.dat" ;
		aph_490_bias:ref = "http://www.uncertweb.org" ;
		aph_490_bias:rel = "uncertainty" ;
		aph_490_bias:units = "m-1" ;
		aph_490_bias:units_nonstandard = "m^-1" ;
		aph_490_bias:wavelength = 490 ;
		aph_490_bias:_Storage = "chunked" ;
		aph_490_bias:_ChunkSizes = 1, 270, 270 ;
		aph_490_bias:_Shuffle = "true" ;
		aph_490_bias:_DeflateLevel = 3 ;
		aph_490_bias:_Endianness = "little" ;
	float aph_490_rmsd(time, lat, lon) ;
		aph_490_rmsd:long_name = "Root-mean-square-difference of phytoplankton absorption coefficient at 490 nm." ;
		aph_490_rmsd:_FillValue = 9.96921e+36f ;
		aph_490_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_rmsd.dat" ;
		aph_490_rmsd:ref = "http://www.uncertweb.org" ;
		aph_490_rmsd:rel = "uncertainty" ;
		aph_490_rmsd:units = "m-1" ;
		aph_490_rmsd:units_nonstandard = "m^-1" ;
		aph_490_rmsd:wavelength = 490 ;
		aph_490_rmsd:_Storage = "chunked" ;
		aph_490_rmsd:_ChunkSizes = 1, 270, 270 ;
		aph_490_rmsd:_Shuffle = "true" ;
		aph_490_rmsd:_DeflateLevel = 3 ;
		aph_490_rmsd:_Endianness = "little" ;
	float aph_510(time, lat, lon) ;
		aph_510:_FillValue = 9.96921e+36f ;
		aph_510:ancillary_variables = "aph_510_rmsd aph_510_bias" ;
		aph_510:grid_mapping = "crs" ;
		aph_510:long_name = "Phytoplankton absorption coefficient at 510 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		aph_510:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		aph_510:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		aph_510:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		aph_510:units = "m-1" ;
		aph_510:units_nonstandard = "m^-1" ;
		aph_510:wavelength = 510 ;
		aph_510:_Storage = "chunked" ;
		aph_510:_ChunkSizes = 1, 270, 270 ;
		aph_510:_Shuffle = "true" ;
		aph_510:_DeflateLevel = 3 ;
		aph_510:_Endianness = "little" ;
	float aph_510_bias(time, lat, lon) ;
		aph_510_bias:long_name = "Bias of phytoplankton absorption coefficient at 510 nm." ;
		aph_510_bias:_FillValue = 9.96921e+36f ;
		aph_510_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_bias.dat" ;
		aph_510_bias:ref = "http://www.uncertweb.org" ;
		aph_510_bias:rel = "uncertainty" ;
		aph_510_bias:units = "m-1" ;
		aph_510_bias:units_nonstandard = "m^-1" ;
		aph_510_bias:wavelength = 510 ;
		aph_510_bias:_Storage = "chunked" ;
		aph_510_bias:_ChunkSizes = 1, 270, 270 ;
		aph_510_bias:_Shuffle = "true" ;
		aph_510_bias:_DeflateLevel = 3 ;
		aph_510_bias:_Endianness = "little" ;
	float aph_510_rmsd(time, lat, lon) ;
		aph_510_rmsd:long_name = "Root-mean-square-difference of phytoplankton absorption coefficient at 510 nm." ;
		aph_510_rmsd:_FillValue = 9.96921e+36f ;
		aph_510_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_rmsd.dat" ;
		aph_510_rmsd:ref = "http://www.uncertweb.org" ;
		aph_510_rmsd:rel = "uncertainty" ;
		aph_510_rmsd:units = "m-1" ;
		aph_510_rmsd:units_nonstandard = "m^-1" ;
		aph_510_rmsd:wavelength = 510 ;
		aph_510_rmsd:_Storage = "chunked" ;
		aph_510_rmsd:_ChunkSizes = 1, 270, 270 ;
		aph_510_rmsd:_Shuffle = "true" ;
		aph_510_rmsd:_DeflateLevel = 3 ;
		aph_510_rmsd:_Endianness = "little" ;
	float aph_560(time, lat, lon) ;
		aph_560:_FillValue = 9.96921e+36f ;
		aph_560:ancillary_variables = "aph_560_rmsd aph_560_bias" ;
		aph_560:grid_mapping = "crs" ;
		aph_560:long_name = "Phytoplankton absorption coefficient at 560 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		aph_560:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		aph_560:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		aph_560:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		aph_560:units = "m-1" ;
		aph_560:units_nonstandard = "m^-1" ;
		aph_560:wavelength = 560 ;
		aph_560:_Storage = "chunked" ;
		aph_560:_ChunkSizes = 1, 270, 270 ;
		aph_560:_Shuffle = "true" ;
		aph_560:_DeflateLevel = 3 ;
		aph_560:_Endianness = "little" ;
	float aph_560_bias(time, lat, lon) ;
		aph_560_bias:long_name = "Bias of phytoplankton absorption coefficient at 560 nm." ;
		aph_560_bias:_FillValue = 9.96921e+36f ;
		aph_560_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_bias.dat" ;
		aph_560_bias:ref = "http://www.uncertweb.org" ;
		aph_560_bias:rel = "uncertainty" ;
		aph_560_bias:units = "m-1" ;
		aph_560_bias:units_nonstandard = "m^-1" ;
		aph_560_bias:wavelength = 560 ;
		aph_560_bias:_Storage = "chunked" ;
		aph_560_bias:_ChunkSizes = 1, 270, 270 ;
		aph_560_bias:_Shuffle = "true" ;
		aph_560_bias:_DeflateLevel = 3 ;
		aph_560_bias:_Endianness = "little" ;
	float aph_560_rmsd(time, lat, lon) ;
		aph_560_rmsd:long_name = "Root-mean-square-difference of phytoplankton absorption coefficient at 560 nm." ;
		aph_560_rmsd:_FillValue = 9.96921e+36f ;
		aph_560_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_rmsd.dat" ;
		aph_560_rmsd:ref = "http://www.uncertweb.org" ;
		aph_560_rmsd:rel = "uncertainty" ;
		aph_560_rmsd:units = "m-1" ;
		aph_560_rmsd:units_nonstandard = "m^-1" ;
		aph_560_rmsd:wavelength = 560 ;
		aph_560_rmsd:_Storage = "chunked" ;
		aph_560_rmsd:_ChunkSizes = 1, 270, 270 ;
		aph_560_rmsd:_Shuffle = "true" ;
		aph_560_rmsd:_DeflateLevel = 3 ;
		aph_560_rmsd:_Endianness = "little" ;
	float aph_665(time, lat, lon) ;
		aph_665:_FillValue = 9.96921e+36f ;
		aph_665:ancillary_variables = "aph_665_rmsd aph_665_bias" ;
		aph_665:grid_mapping = "crs" ;
		aph_665:long_name = "Phytoplankton absorption coefficient at 665 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		aph_665:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		aph_665:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0063" ;
		aph_665:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		aph_665:units = "m-1" ;
		aph_665:units_nonstandard = "m^-1" ;
		aph_665:wavelength = 665 ;
		aph_665:_Storage = "chunked" ;
		aph_665:_ChunkSizes = 1, 270, 270 ;
		aph_665:_Shuffle = "true" ;
		aph_665:_DeflateLevel = 3 ;
		aph_665:_Endianness = "little" ;
	float aph_665_bias(time, lat, lon) ;
		aph_665_bias:long_name = "Bias of phytoplankton absorption coefficient at 665 nm." ;
		aph_665_bias:_FillValue = 9.96921e+36f ;
		aph_665_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_bias.dat" ;
		aph_665_bias:ref = "http://www.uncertweb.org" ;
		aph_665_bias:rel = "uncertainty" ;
		aph_665_bias:units = "m-1" ;
		aph_665_bias:units_nonstandard = "m^-1" ;
		aph_665_bias:wavelength = 665 ;
		aph_665_bias:_Storage = "chunked" ;
		aph_665_bias:_ChunkSizes = 1, 270, 270 ;
		aph_665_bias:_Shuffle = "true" ;
		aph_665_bias:_DeflateLevel = 3 ;
		aph_665_bias:_Endianness = "little" ;
	float aph_665_rmsd(time, lat, lon) ;
		aph_665_rmsd:long_name = "Root-mean-square-difference of phytoplankton absorption coefficient at 665 nm." ;
		aph_665_rmsd:_FillValue = 9.96921e+36f ;
		aph_665_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/aph/cci_iop_aph_rmsd.dat" ;
		aph_665_rmsd:ref = "http://www.uncertweb.org" ;
		aph_665_rmsd:rel = "uncertainty" ;
		aph_665_rmsd:units = "m-1" ;
		aph_665_rmsd:units_nonstandard = "m^-1" ;
		aph_665_rmsd:wavelength = 665 ;
		aph_665_rmsd:_Storage = "chunked" ;
		aph_665_rmsd:_ChunkSizes = 1, 270, 270 ;
		aph_665_rmsd:_Shuffle = "true" ;
		aph_665_rmsd:_DeflateLevel = 3 ;
		aph_665_rmsd:_Endianness = "little" ;
	float atot_412(time, lat, lon) ;
		atot_412:_FillValue = 9.96921e+36f ;
		atot_412:long_name = "Total absorption coefficient at 412 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		atot_412:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		atot_412:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0062" ;
		atot_412:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		atot_412:units = "m-1" ;
		atot_412:units_nonstandard = "m^-1" ;
		atot_412:wavelength = 412 ;
		atot_412:_Storage = "chunked" ;
		atot_412:_ChunkSizes = 1, 270, 270 ;
		atot_412:_Shuffle = "true" ;
		atot_412:_DeflateLevel = 3 ;
		atot_412:_Endianness = "little" ;
	float atot_443(time, lat, lon) ;
		atot_443:_FillValue = 9.96921e+36f ;
		atot_443:long_name = "Total absorption coefficient at 443 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		atot_443:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		atot_443:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0062" ;
		atot_443:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		atot_443:units = "m-1" ;
		atot_443:units_nonstandard = "m^-1" ;
		atot_443:wavelength = 443 ;
		atot_443:_Storage = "chunked" ;
		atot_443:_ChunkSizes = 1, 270, 270 ;
		atot_443:_Shuffle = "true" ;
		atot_443:_DeflateLevel = 3 ;
		atot_443:_Endianness = "little" ;
	float atot_490(time, lat, lon) ;
		atot_490:_FillValue = 9.96921e+36f ;
		atot_490:long_name = "Total absorption coefficient at 490 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		atot_490:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		atot_490:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0062" ;
		atot_490:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		atot_490:units = "m-1" ;
		atot_490:units_nonstandard = "m^-1" ;
		atot_490:wavelength = 490 ;
		atot_490:_Storage = "chunked" ;
		atot_490:_ChunkSizes = 1, 270, 270 ;
		atot_490:_Shuffle = "true" ;
		atot_490:_DeflateLevel = 3 ;
		atot_490:_Endianness = "little" ;
	float atot_510(time, lat, lon) ;
		atot_510:_FillValue = 9.96921e+36f ;
		atot_510:long_name = "Total absorption coefficient at 510 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		atot_510:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		atot_510:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0062" ;
		atot_510:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		atot_510:units = "m-1" ;
		atot_510:units_nonstandard = "m^-1" ;
		atot_510:wavelength = 510 ;
		atot_510:_Storage = "chunked" ;
		atot_510:_ChunkSizes = 1, 270, 270 ;
		atot_510:_Shuffle = "true" ;
		atot_510:_DeflateLevel = 3 ;
		atot_510:_Endianness = "little" ;
	float atot_560(time, lat, lon) ;
		atot_560:_FillValue = 9.96921e+36f ;
		atot_560:long_name = "Total absorption coefficient at 560 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		atot_560:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		atot_560:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0062" ;
		atot_560:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		atot_560:units = "m-1" ;
		atot_560:units_nonstandard = "m^-1" ;
		atot_560:wavelength = 560 ;
		atot_560:_Storage = "chunked" ;
		atot_560:_ChunkSizes = 1, 270, 270 ;
		atot_560:_Shuffle = "true" ;
		atot_560:_DeflateLevel = 3 ;
		atot_560:_Endianness = "little" ;
	float atot_665(time, lat, lon) ;
		atot_665:_FillValue = 9.96921e+36f ;
		atot_665:long_name = "Total absorption coefficient at 665 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		atot_665:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		atot_665:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0062" ;
		atot_665:standard_name = "volume_absorption_coefficient_of_radiative_flux_in_sea_water" ;
		atot_665:units = "m-1" ;
		atot_665:units_nonstandard = "m^-1" ;
		atot_665:wavelength = 665 ;
		atot_665:_Storage = "chunked" ;
		atot_665:_ChunkSizes = 1, 270, 270 ;
		atot_665:_Shuffle = "true" ;
		atot_665:_DeflateLevel = 3 ;
		atot_665:_Endianness = "little" ;
	float bbp_412(time, lat, lon) ;
		bbp_412:_FillValue = 9.96921e+36f ;
		bbp_412:long_name = "Particulate backscattering coefficient for dissolved and detrital material at 412 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		bbp_412:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		bbp_412:parameter_vocab_uri = "http://vocab.nerc.ac.uk/collection/P04/current/" ;
		bbp_412:standard_name = "volume_backwards_scattering_coefficient_of_radiative_flux_in_sea_water" ;
		bbp_412:units = "m-1" ;
		bbp_412:units_nonstandard = "m^-1" ;
		bbp_412:wavelength = 412 ;
		bbp_412:_Storage = "chunked" ;
		bbp_412:_ChunkSizes = 1, 270, 270 ;
		bbp_412:_Shuffle = "true" ;
		bbp_412:_DeflateLevel = 3 ;
		bbp_412:_Endianness = "little" ;
	float bbp_443(time, lat, lon) ;
		bbp_443:_FillValue = 9.96921e+36f ;
		bbp_443:long_name = "Particulate backscattering coefficient for dissolved and detrital material at 443 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		bbp_443:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		bbp_443:parameter_vocab_uri = "http://vocab.nerc.ac.uk/collection/P04/current/" ;
		bbp_443:standard_name = "volume_backwards_scattering_coefficient_of_radiative_flux_in_sea_water" ;
		bbp_443:units = "m-1" ;
		bbp_443:units_nonstandard = "m^-1" ;
		bbp_443:wavelength = 443 ;
		bbp_443:_Storage = "chunked" ;
		bbp_443:_ChunkSizes = 1, 270, 270 ;
		bbp_443:_Shuffle = "true" ;
		bbp_443:_DeflateLevel = 3 ;
		bbp_443:_Endianness = "little" ;
	float bbp_490(time, lat, lon) ;
		bbp_490:_FillValue = 9.96921e+36f ;
		bbp_490:long_name = "Particulate backscattering coefficient for dissolved and detrital material at 490 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		bbp_490:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		bbp_490:parameter_vocab_uri = "http://vocab.nerc.ac.uk/collection/P04/current/" ;
		bbp_490:standard_name = "volume_backwards_scattering_coefficient_of_radiative_flux_in_sea_water" ;
		bbp_490:units = "m-1" ;
		bbp_490:units_nonstandard = "m^-1" ;
		bbp_490:wavelength = 490 ;
		bbp_490:_Storage = "chunked" ;
		bbp_490:_ChunkSizes = 1, 270, 270 ;
		bbp_490:_Shuffle = "true" ;
		bbp_490:_DeflateLevel = 3 ;
		bbp_490:_Endianness = "little" ;
	float bbp_510(time, lat, lon) ;
		bbp_510:_FillValue = 9.96921e+36f ;
		bbp_510:long_name = "Particulate backscattering coefficient for dissolved and detrital material at 510 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		bbp_510:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		bbp_510:parameter_vocab_uri = "http://vocab.nerc.ac.uk/collection/P04/current/" ;
		bbp_510:standard_name = "volume_backwards_scattering_coefficient_of_radiative_flux_in_sea_water" ;
		bbp_510:units = "m-1" ;
		bbp_510:units_nonstandard = "m^-1" ;
		bbp_510:wavelength = 510 ;
		bbp_510:_Storage = "chunked" ;
		bbp_510:_ChunkSizes = 1, 270, 270 ;
		bbp_510:_Shuffle = "true" ;
		bbp_510:_DeflateLevel = 3 ;
		bbp_510:_Endianness = "little" ;
	float bbp_560(time, lat, lon) ;
		bbp_560:_FillValue = 9.96921e+36f ;
		bbp_560:long_name = "Particulate backscattering coefficient for dissolved and detrital material at 560 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		bbp_560:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		bbp_560:parameter_vocab_uri = "http://vocab.nerc.ac.uk/collection/P04/current/" ;
		bbp_560:standard_name = "volume_backwards_scattering_coefficient_of_radiative_flux_in_sea_water" ;
		bbp_560:units = "m-1" ;
		bbp_560:units_nonstandard = "m^-1" ;
		bbp_560:wavelength = 560 ;
		bbp_560:_Storage = "chunked" ;
		bbp_560:_ChunkSizes = 1, 270, 270 ;
		bbp_560:_Shuffle = "true" ;
		bbp_560:_DeflateLevel = 3 ;
		bbp_560:_Endianness = "little" ;
	float bbp_665(time, lat, lon) ;
		bbp_665:_FillValue = 9.96921e+36f ;
		bbp_665:long_name = "Particulate backscattering coefficient for dissolved and detrital material at 665 nm derived using the QAA model V6 (Lee et al 2014) as parameterised within SeaDAS." ;
		bbp_665:paper_ref = "Lee, Z., et al. Update of the Quasi-Analytical Algorithm (QAA_v6) [R/OL]. International Ocean Color Group Software Report [2013-04-03]. http://www.ioccg.org/groups/Software-OCA/OAA_5.2014." ;
		bbp_665:parameter_vocab_uri = "http://vocab.nerc.ac.uk/collection/P04/current/" ;
		bbp_665:standard_name = "volume_backwards_scattering_coefficient_of_radiative_flux_in_sea_water" ;
		bbp_665:units = "m-1" ;
		bbp_665:units_nonstandard = "m^-1" ;
		bbp_665:wavelength = 665 ;
		bbp_665:_Storage = "chunked" ;
		bbp_665:_ChunkSizes = 1, 270, 270 ;
		bbp_665:_Shuffle = "true" ;
		bbp_665:_DeflateLevel = 3 ;
		bbp_665:_Endianness = "little" ;
	float chlor_a(time, lat, lon) ;
		chlor_a:_FillValue = 9.96921e+36f ;
		chlor_a:ancillary_variables = "chlor_a_log10_rmsd chlor_a_log10_bias" ;
		chlor_a:long_name = "Chlorophyll-a concentration in seawater (not log-transformed), generated by as a blended combination of OCI, OCI2, OC2 and OCx algorithms, depending on water class memberships" ;
		chlor_a:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P011/current/CHLTVOLU" ;
		chlor_a:standard_name = "mass_concentration_of_chlorophyll_a_in_sea_water" ;
		chlor_a:units = "milligram m-3" ;
		chlor_a:units_nonstandard = "mg m^-3" ;
		chlor_a:_Storage = "chunked" ;
		chlor_a:_ChunkSizes = 1, 270, 270 ;
		chlor_a:_Shuffle = "true" ;
		chlor_a:_DeflateLevel = 3 ;
		chlor_a:_Endianness = "little" ;
	float chlor_a_log10_bias(time, lat, lon) ;
		chlor_a_log10_bias:long_name = "Bias of log10-transformed chlorophyll-a concentration in seawater." ;
		chlor_a_log10_bias:_FillValue = 9.96921e+36f ;
		chlor_a_log10_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/chlor_a/cci_chla_bias.dat" ;
		chlor_a_log10_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		chlor_a_log10_bias:rel = "uncertainty" ;
		chlor_a_log10_bias:_Storage = "chunked" ;
		chlor_a_log10_bias:_ChunkSizes = 1, 270, 270 ;
		chlor_a_log10_bias:_Shuffle = "true" ;
		chlor_a_log10_bias:_DeflateLevel = 3 ;
		chlor_a_log10_bias:_Endianness = "little" ;
	float chlor_a_log10_rmsd(time, lat, lon) ;
		chlor_a_log10_rmsd:long_name = "Root-mean-square-difference of log10-transformed chlorophyll-a concentration in seawater." ;
		chlor_a_log10_rmsd:_FillValue = 9.96921e+36f ;
		chlor_a_log10_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/chlor_a/cci_chla_rmsd.dat" ;
		chlor_a_log10_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		chlor_a_log10_rmsd:rel = "uncertainty" ;
		chlor_a_log10_rmsd:_Storage = "chunked" ;
		chlor_a_log10_rmsd:_ChunkSizes = 1, 270, 270 ;
		chlor_a_log10_rmsd:_Shuffle = "true" ;
		chlor_a_log10_rmsd:_DeflateLevel = 3 ;
		chlor_a_log10_rmsd:_Endianness = "little" ;
	float kd_490(time, lat, lon) ;
		kd_490:_FillValue = 9.96921e+36f ;
		kd_490:ancillary_variables = "kd_490_rmsd kd_490_bias" ;
		kd_490:long_name = "Downwelling attenuation coefficient at 490nm, derived using Lee 2005 equation and bbw from Zhang 2009 (following the SeaDAS Kd_lee algorithm)" ;
		kd_490:parameter_vocab_uri = "http://vocab.ndg.nerc.ac.uk/term/P071/19/CFSN0064" ;
		kd_490:standard_name = "volume_attenuation_coefficient_of_downwelling_radiative_flux_in_sea_water" ;
		kd_490:units = "m-1" ;
		kd_490:units_nonstandard = "m^-1" ;
		kd_490:wavelength = 490 ;
		kd_490:_Storage = "chunked" ;
		kd_490:_ChunkSizes = 1, 270, 270 ;
		kd_490:_Shuffle = "true" ;
		kd_490:_DeflateLevel = 3 ;
		kd_490:_Endianness = "little" ;
	float kd_490_bias(time, lat, lon) ;
		kd_490_bias:long_name = "Bias of downwelling attenuation coefficient at 490 nm derived using Lee 2005 equation and bbw from Zhang 2009" ;
		kd_490_bias:_FillValue = 9.96921e+36f ;
		kd_490_bias:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/kd/cci_kd_bias.dat" ;
		kd_490_bias:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		kd_490_bias:rel = "uncertainty" ;
		kd_490_bias:units = "m-1" ;
		kd_490_bias:units_nonstandard = "m^-1" ;
		kd_490_bias:wavelength = 490 ;
		kd_490_bias:_Storage = "chunked" ;
		kd_490_bias:_ChunkSizes = 1, 270, 270 ;
		kd_490_bias:_Shuffle = "true" ;
		kd_490_bias:_DeflateLevel = 3 ;
		kd_490_bias:_Endianness = "little" ;
	float kd_490_rmsd(time, lat, lon) ;
		kd_490_rmsd:long_name = "Root-mean-square-difference of downwelling attenuation coefficient at 490 nm derived using Lee 2005 equation and bbw from Zhang 2009" ;
		kd_490_rmsd:_FillValue = 9.96921e+36f ;
		kd_490_rmsd:comment = "Uncertainty lookups derived from file: /data/datasets/CCI/v6.0-production/stage09b-uncertainty_tables/kd/cci_kd_rmsd.dat" ;
		kd_490_rmsd:ref = "http://www.esa-oceancolour-cci.org/?q=webfm_send/581" ;
		kd_490_rmsd:rel = "uncertainty" ;
		kd_490_rmsd:units = "m-1" ;
		kd_490_rmsd:units_nonstandard = "m^-1" ;
		kd_490_rmsd:wavelength = 490 ;
		kd_490_rmsd:_Storage = "chunked" ;
		kd_490_rmsd:_ChunkSizes = 1, 270, 270 ;
		kd_490_rmsd:_Shuffle = "true" ;
		kd_490_rmsd:_DeflateLevel = 3 ;
		kd_490_rmsd:_Endianness = "little" ;
	double lat(lat) ;
		lat:units = "degrees_north" ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:valid_min = -89.9791666666667 ;
		lat:valid_max = 89.9791666666667 ;
		lat:axis = "Y" ;
		lat:_Storage = "chunked" ;
		lat:_ChunkSizes = 270 ;
		lat:_Shuffle = "true" ;
		lat:_DeflateLevel = 3 ;
		lat:_Endianness = "little" ;
	double lon(lon) ;
		lon:units = "degrees_east" ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:valid_min = -179.979166666667 ;
		lon:valid_max = 179.979166666667 ;
		lon:axis = "X" ;
		lon:_Storage = "chunked" ;
		lon:_ChunkSizes = 270 ;
		lon:_Shuffle = "true" ;
		lon:_DeflateLevel = 3 ;
		lon:_Endianness = "little" ;
	int time(time) ;
		time:axis = "T" ;
		time:standard_name = "time" ;
		time:units = "days since 1970-01-01 00:00:00" ;
		time:_Storage = "chunked" ;
		time:_ChunkSizes = 1 ;
		time:_Shuffle = "true" ;
		time:_DeflateLevel = 3 ;
		time:_Endianness = "little" ;
	float water_class1(time, lat, lon) ;
		water_class1:_FillValue = 9.96921e+36f ;
		water_class1:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class1:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class1:long_name = "Mean of normalised water class 1 membership over the compositing period" ;
		water_class1:_Storage = "chunked" ;
		water_class1:_ChunkSizes = 1, 270, 270 ;
		water_class1:_Shuffle = "true" ;
		water_class1:_DeflateLevel = 3 ;
		water_class1:_Endianness = "little" ;
	float water_class10(time, lat, lon) ;
		water_class10:_FillValue = 9.96921e+36f ;
		water_class10:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class10:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class10:long_name = "Mean of normalised water class 10 membership over the compositing period" ;
		water_class10:_Storage = "chunked" ;
		water_class10:_ChunkSizes = 1, 270, 270 ;
		water_class10:_Shuffle = "true" ;
		water_class10:_DeflateLevel = 3 ;
		water_class10:_Endianness = "little" ;
	float water_class11(time, lat, lon) ;
		water_class11:_FillValue = 9.96921e+36f ;
		water_class11:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class11:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class11:long_name = "Mean of normalised water class 11 membership over the compositing period" ;
		water_class11:_Storage = "chunked" ;
		water_class11:_ChunkSizes = 1, 270, 270 ;
		water_class11:_Shuffle = "true" ;
		water_class11:_DeflateLevel = 3 ;
		water_class11:_Endianness = "little" ;
	float water_class12(time, lat, lon) ;
		water_class12:_FillValue = 9.96921e+36f ;
		water_class12:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class12:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class12:long_name = "Mean of normalised water class 12 membership over the compositing period" ;
		water_class12:_Storage = "chunked" ;
		water_class12:_ChunkSizes = 1, 270, 270 ;
		water_class12:_Shuffle = "true" ;
		water_class12:_DeflateLevel = 3 ;
		water_class12:_Endianness = "little" ;
	float water_class13(time, lat, lon) ;
		water_class13:_FillValue = 9.96921e+36f ;
		water_class13:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class13:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class13:long_name = "Mean of normalised water class 13 membership over the compositing period" ;
		water_class13:_Storage = "chunked" ;
		water_class13:_ChunkSizes = 1, 270, 270 ;
		water_class13:_Shuffle = "true" ;
		water_class13:_DeflateLevel = 3 ;
		water_class13:_Endianness = "little" ;
	float water_class14(time, lat, lon) ;
		water_class14:_FillValue = 9.96921e+36f ;
		water_class14:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class14:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class14:long_name = "Mean of normalised water class 14 membership over the compositing period" ;
		water_class14:_Storage = "chunked" ;
		water_class14:_ChunkSizes = 1, 270, 270 ;
		water_class14:_Shuffle = "true" ;
		water_class14:_DeflateLevel = 3 ;
		water_class14:_Endianness = "little" ;
	float water_class2(time, lat, lon) ;
		water_class2:_FillValue = 9.96921e+36f ;
		water_class2:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class2:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class2:long_name = "Mean of normalised water class 2 membership over the compositing period" ;
		water_class2:_Storage = "chunked" ;
		water_class2:_ChunkSizes = 1, 270, 270 ;
		water_class2:_Shuffle = "true" ;
		water_class2:_DeflateLevel = 3 ;
		water_class2:_Endianness = "little" ;
	float water_class3(time, lat, lon) ;
		water_class3:_FillValue = 9.96921e+36f ;
		water_class3:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class3:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class3:long_name = "Mean of normalised water class 3 membership over the compositing period" ;
		water_class3:_Storage = "chunked" ;
		water_class3:_ChunkSizes = 1, 270, 270 ;
		water_class3:_Shuffle = "true" ;
		water_class3:_DeflateLevel = 3 ;
		water_class3:_Endianness = "little" ;
	float water_class4(time, lat, lon) ;
		water_class4:_FillValue = 9.96921e+36f ;
		water_class4:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class4:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class4:long_name = "Mean of normalised water class 4 membership over the compositing period" ;
		water_class4:_Storage = "chunked" ;
		water_class4:_ChunkSizes = 1, 270, 270 ;
		water_class4:_Shuffle = "true" ;
		water_class4:_DeflateLevel = 3 ;
		water_class4:_Endianness = "little" ;
	float water_class5(time, lat, lon) ;
		water_class5:_FillValue = 9.96921e+36f ;
		water_class5:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class5:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class5:long_name = "Mean of normalised water class 5 membership over the compositing period" ;
		water_class5:_Storage = "chunked" ;
		water_class5:_ChunkSizes = 1, 270, 270 ;
		water_class5:_Shuffle = "true" ;
		water_class5:_DeflateLevel = 3 ;
		water_class5:_Endianness = "little" ;
	float water_class6(time, lat, lon) ;
		water_class6:_FillValue = 9.96921e+36f ;
		water_class6:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class6:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class6:long_name = "Mean of normalised water class 6 membership over the compositing period" ;
		water_class6:_Storage = "chunked" ;
		water_class6:_ChunkSizes = 1, 270, 270 ;
		water_class6:_Shuffle = "true" ;
		water_class6:_DeflateLevel = 3 ;
		water_class6:_Endianness = "little" ;
	float water_class7(time, lat, lon) ;
		water_class7:_FillValue = 9.96921e+36f ;
		water_class7:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class7:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class7:long_name = "Mean of normalised water class 7 membership over the compositing period" ;
		water_class7:_Storage = "chunked" ;
		water_class7:_ChunkSizes = 1, 270, 270 ;
		water_class7:_Shuffle = "true" ;
		water_class7:_DeflateLevel = 3 ;
		water_class7:_Endianness = "little" ;
	float water_class8(time, lat, lon) ;
		water_class8:_FillValue = 9.96921e+36f ;
		water_class8:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class8:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class8:long_name = "Mean of normalised water class 8 membership over the compositing period" ;
		water_class8:_Storage = "chunked" ;
		water_class8:_ChunkSizes = 1, 270, 270 ;
		water_class8:_Shuffle = "true" ;
		water_class8:_DeflateLevel = 3 ;
		water_class8:_Endianness = "little" ;
	float water_class9(time, lat, lon) ;
		water_class9:_FillValue = 9.96921e+36f ;
		water_class9:paper_ref = "Thomas Jackson, Shubha Sathyendranath, Frederic Melin, (2017) An improved optical classification scheme for the Ocean Colour Essential Climate Variable and its applications, Remote Sensing of Environment, Available online 5 April 2017, ISSN 0034-4257, http://doi.org/10.1016/j.rse.2017.03.036." ;
		water_class9:ref = "http://dx.doi.org/10.1016/j.rse.2009.07.016" ;
		water_class9:long_name = "Mean of normalised water class 9 membership over the compositing period" ;
		water_class9:_Storage = "chunked" ;
		water_class9:_ChunkSizes = 1, 270, 270 ;
		water_class9:_Shuffle = "true" ;
		water_class9:_DeflateLevel = 3 ;
		water_class9:_Endianness = "little" ;
	int crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:_Storage = "contiguous" ;
		crs:_Endianness = "little" ;
	float MERIS_nobs_sum(time, lat, lon) ;
		MERIS_nobs_sum:_FillValue = 0.f ;
		MERIS_nobs_sum:long_name = "Count of the number of observations from the MERIS sensor contributing to this bin cell" ;
		MERIS_nobs_sum:number_of_files_composited = 31 ;
		MERIS_nobs_sum:_Storage = "chunked" ;
		MERIS_nobs_sum:_ChunkSizes = 1, 270, 270 ;
		MERIS_nobs_sum:_Shuffle = "true" ;
		MERIS_nobs_sum:_DeflateLevel = 3 ;
		MERIS_nobs_sum:_Endianness = "little" ;
	float MODISA_nobs_sum(time, lat, lon) ;
		MODISA_nobs_sum:_FillValue = 0.f ;
		MODISA_nobs_sum:long_name = "Count of the number of observations from the MODIS (Aqua) sensor contributing to this bin cell" ;
		MODISA_nobs_sum:number_of_files_composited = 31 ;
		MODISA_nobs_sum:_Storage = "chunked" ;
		MODISA_nobs_sum:_ChunkSizes = 1, 270, 270 ;
		MODISA_nobs_sum:_Shuffle = "true" ;
		MODISA_nobs_sum:_DeflateLevel = 3 ;
		MODISA_nobs_sum:_Endianness = "little" ;
	float OLCI-A_nobs_sum(time, lat, lon) ;
		OLCI-A_nobs_sum:_FillValue = 0.f ;
		OLCI-A_nobs_sum:long_name = "Count of the number of observations from the OLCI (Sentinel-3a) sensor contributing to this bin cell" ;
		OLCI-A_nobs_sum:number_of_files_composited = 31 ;
		OLCI-A_nobs_sum:_Storage = "chunked" ;
		OLCI-A_nobs_sum:_ChunkSizes = 1, 270, 270 ;
		OLCI-A_nobs_sum:_Shuffle = "true" ;
		OLCI-A_nobs_sum:_DeflateLevel = 3 ;
		OLCI-A_nobs_sum:_Endianness = "little" ;
	float OLCI-B_nobs_sum(time, lat, lon) ;
		OLCI-B_nobs_sum:_FillValue = 0.f ;
		OLCI-B_nobs_sum:long_name = "Count of the number of observations from the OLCI (Sentinel-3b) sensor contributing to this bin cell" ;
		OLCI-B_nobs_sum:number_of_files_composited = 31 ;
		OLCI-B_nobs_sum:_Storage = "chunked" ;
		OLCI-B_nobs_sum:_ChunkSizes = 1, 270, 270 ;
		OLCI-B_nobs_sum:_Shuffle = "true" ;
		OLCI-B_nobs_sum:_DeflateLevel = 3 ;
		OLCI-B_nobs_sum:_Endianness = "little" ;
	float SeaWiFS_nobs_sum(time, lat, lon) ;
		SeaWiFS_nobs_sum:_FillValue = 0.f ;
		SeaWiFS_nobs_sum:long_name = "Count of the number of observations from the SeaWiFS (GAC and LAC) sensor contributing to this bin cell" ;
		SeaWiFS_nobs_sum:number_of_files_composited = 31 ;
		SeaWiFS_nobs_sum:_Storage = "chunked" ;
		SeaWiFS_nobs_sum:_ChunkSizes = 1, 270, 270 ;
		SeaWiFS_nobs_sum:_Shuffle = "true" ;
		SeaWiFS_nobs_sum:_DeflateLevel = 3 ;
		SeaWiFS_nobs_sum:_Endianness = "little" ;
	float VIIRS_nobs_sum(time, lat, lon) ;
		VIIRS_nobs_sum:_FillValue = 0.f ;
		VIIRS_nobs_sum:long_name = "Count of the number of observations from the VIIRS sensor contributing to this bin cell" ;
		VIIRS_nobs_sum:number_of_files_composited = 31 ;
		VIIRS_nobs_sum:_Storage = "chunked" ;
		VIIRS_nobs_sum:_ChunkSizes = 1, 270, 270 ;
		VIIRS_nobs_sum:_Shuffle = "true" ;
		VIIRS_nobs_sum:_DeflateLevel = 3 ;
		VIIRS_nobs_sum:_Endianness = "little" ;
	float total_nobs_sum(time, lat, lon) ;
		total_nobs_sum:_FillValue = 0.f ;
		total_nobs_sum:long_name = "Count of the total number of observations contributing to this bin cell" ;
		total_nobs_sum:number_of_files_composited = 31 ;
		total_nobs_sum:_Storage = "chunked" ;
		total_nobs_sum:_ChunkSizes = 1, 270, 270 ;
		total_nobs_sum:_Shuffle = "true" ;
		total_nobs_sum:_DeflateLevel = 3 ;
		total_nobs_sum:_Endianness = "little" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:cdm_data_type = "Grid" ;
		:comment = "See summary attribute" ;
		:creator_email = "help@esa-oceancolour-cci.org" ;
		:creator_name = "Plymouth Marine Laboratory" ;
		:creator_url = "http://esa-oceancolour-cci.org" ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lat_resolution = ".04166666666666666666" ;
		:geospatial_lat_units = "decimal degrees north" ;
		:geospatial_lon_max = 180.f ;
		:geospatial_lon_min = -180.f ;
		:geospatial_lon_resolution = ".04166666666666666666" ;
		:geospatial_lon_units = "decimal degrees east" ;
		:geospatial_vertical_max = 0.f ;
		:geospatial_vertical_min = 0.f ;
		:git_commit_hash = "4db7bf1d93d4acce920d50186c81b2052007f64a" ;
		:institution = "Plymouth Marine Laboratory" ;
		:keywords = "satellite,observation,ocean,ocean colour" ;
		:keywords_vocabulary = "none" ;
		:license = "ESA CCI Data Policy: free and open access.  When referencing, please use: Ocean Colour Climate Change Initiative dataset, Version <Version Number>, European Space Agency, available online at http://www.esa-oceancolour-cci.org.  We would also appreciate being notified of publications so that we can list them on the project website at http://www.esa-oceancolour-cci.org/?q=publications" ;
		:naming_authority = "uk.ac.pml" ;
		:number_of_bands_used_to_classify = "4" ;
		:number_of_optical_water_types = "14" ;
		:platform = "Orbview-2,Aqua,Envisat,Suomi-NPP, Sentinel-3a, Sentinel-3b" ;
		:processing_level = "Level-3" ;
		:product_version = "6.0" ;
		:project = "Climate Change Initiative - European Space Agency" ;
		:references = "http://www.esa-oceancolour-cci.org/" ;
		:sensor = "SeaWiFS,MODIS,MERIS,VIIRS,OLCI" ;
		:sensors_present = " SeaWiFS" ;
		:spatial_resolution = "4km nominal at equator" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Conventions Version 1.7" ;
		:title = "ESA CCI Ocean Colour Product" ;
		:NCO = "netCDF Operators version 4.7.5 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
		:number_of_files_composited = 31 ;
		:history = "Source data were: ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000101-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000102-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000103-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000104-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000105-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000106-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000107-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000108-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000109-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000110-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000111-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000112-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000113-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000114-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000115-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000116-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000117-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000118-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000119-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000120-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000121-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000122-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000123-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000124-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000125-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000126-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000127-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000128-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000129-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000130-fv6.0.nc, ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1D_DAILY_4km_GEO_PML_OCx_QAA-20000131-fv6.0.nc; netcdf_compositor_cci composites  Rrs_412, Rrs_412_bias, Rrs_443, Rrs_443_bias, Rrs_490, Rrs_490_bias, Rrs_510, Rrs_510_bias, Rrs_560, Rrs_560_bias, Rrs_665, Rrs_665_bias, adg_412, adg_412_bias, adg_443, adg_443_bias, adg_490, adg_490_bias, adg_510, adg_510_bias, adg_560, adg_560_bias, adg_665, adg_665_bias, aph_412, aph_412_bias, aph_443, aph_443_bias, aph_490, aph_490_bias, aph_510, aph_510_bias, aph_560, aph_560_bias, aph_665, aph_665_bias, atot_412, atot_443, atot_490, atot_510, atot_560, atot_665, bbp_412, bbp_443, bbp_490, bbp_510, bbp_560, bbp_665, chlor_a, chlor_a_log10_bias, kd_490, kd_490_bias, water_class1, water_class10, water_class11, water_class12, water_class13, water_class14, water_class2, water_class3, water_class4, water_class5, water_class6, water_class7, water_class8, water_class9 with --mean,  Rrs_412_rmsd, Rrs_443_rmsd, Rrs_490_rmsd, Rrs_510_rmsd, Rrs_560_rmsd, Rrs_665_rmsd, adg_412_rmsd, adg_443_rmsd, adg_490_rmsd, adg_510_rmsd, adg_560_rmsd, adg_665_rmsd, aph_412_rmsd, aph_443_rmsd, aph_490_rmsd, aph_510_rmsd, aph_560_rmsd, aph_665_rmsd, chlor_a_log10_rmsd, kd_490_rmsd with --root-mean-square, and  MERIS_nobs, MODISA_nobs, OLCI-A_nobs, OLCI-B_nobs, SeaWiFS_nobs, VIIRS_nobs, total_nobs - with --total" ;
		:id = "ESACCI-OC-L3S-OC_PRODUCTS-MERGED-1M_MONTHLY_4km_GEO_PML_OCx_QAA-200001-fv6.0.nc" ;
		:creation_date = "Mon Aug 15 12:20:17 2022" ;
		:date_created = "Mon Aug 15 12:20:17 2022" ;
		:time_coverage_resolution = "P1M" ;
		:time_coverage_duration = "P1M" ;
		:start_date = "01-JAN-2000 00:00:00.000000" ;
		:stop_date = "31-JAN-2000 23:59:00.000000" ;
		:time_coverage_start = "200001010000Z" ;
		:time_coverage_end = "200001312359Z" ;
		:source = "NASA SeaWiFS  L1A and L2 R2018.0 LAC and GAC, MODIS-Aqua L1A and L2 R2018.0, MERIS L1B 4th reprocessing inc OCL corrections, NASA VIIRS L1A and L2 R2018.0, OLCI L1B" ;
		:summary = "Data products generated by the Ocean Colour component of the European Space Agency Climate Change Initiative project. These files are monthly composites of merged sensor (MERIS, MODIS Aqua, SeaWiFS LAC & GAC, VIIRS, OLCI) products.  MODIS Aqua and SeaWiFS were band-shifted and bias-corrected to MERIS bands and values using a temporally and spatially varying scheme based on the overlap years of 2003-2007.  VIIRS was band-shifted and bias-corrected in a second stage against the MODIS Rrs that had already been corrected to MERIS levels, for the overlap period 2012-2014; at the third stage Sentinel-3A OLCI was bias corrected against already corrected MODIS, for overlap period 2016-07-01 to 2019-06-30;  at the fourth stage Sentinel-3B OLCI was bias corrected against already corrected Sentinel-3A OLCI, for overlap period 2018-07-01 to 2021-06-30.  VIIRS, MODIS, SeaWiFS and MERIS Rrs were derived from a combination of NASA\'s l2gen (for basic sensor geometry corrections, etc) and HYGEOS POLYMER (for atmospheric correction). OLCI Rrs were sourced at L1b (already geometrically corrected) and processed with POLYMER.  The Rrs were binned to a sinusoidal 4km level-3 grid, and later to 4km geographic projection, by Brockmann Consult\'s SNAP.  Derived products were generally computed with the standard algorithms through SeaDAS.  QAA IOPs were derived using the standard SeaDAS algorithm but with a modified backscattering table to match that used in the bandshifting.  The final chlorophyll is a combination of OCI, OCI2, OC2 and OCx, depending on the water class memberships.  Uncertainty estimates were added using the fuzzy water classifier and uncertainty estimation algorithm of Tim Moore as documented in Jackson et al (2017). and updated according to Jackson et al. (in prep)." ;
		:tracking_id = "8d3e6320-4159-4058-87df-ede447dfb6b0" ;
		:_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.20" ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 0 ;
		:_Format = "netCDF-4 classic model" ;
}
