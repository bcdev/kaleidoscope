netcdf Ford_et_al_UExP-FNN-U_physics_carbonatesystem_ESASCOPE_v5 {
dimensions:
	longitude = 360 ;
	latitude = 180 ;
	time = 468 ;
variables:
	float fco2(longitude, latitude, time) ;
		fco2:units = "uatm" ;
		fco2:long_name = "Fugacity of CO2 in seawater" ;
		fco2:comment = "" ;
		fco2:date_variable = "28/02/2025 17:28" ;
		fco2:predictor_parameters = "[\'CCI_SST_analysed_sst\', \'NOAA_ERSL_xCO2\', \'CCI_SSS_sss_CMEMS_so\', \'CMEMS_mlotst\', \'CCI_SST_analysed_sst_anom\', \'NOAA_ERSL_xCO2_anom\', \'CCI_SSS_sss_CMEMS_so_anom\', \'CMEMS_mlotst_anom\']" ;
		fco2:ensemble_size = "10" ;
		fco2:province_variable = "prov_smoothed" ;
		fco2:_Storage = "contiguous" ;
		fco2:_Endianness = "little" ;
	float fco2_net_unc(longitude, latitude, time) ;
		fco2_net_unc:units = "uatm" ;
		fco2_net_unc:long_name = "Fugacity of CO2 in seawater network uncertainty" ;
		fco2_net_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		fco2_net_unc:date_variable = "28/02/2025 17:28" ;
		fco2_net_unc:_Storage = "contiguous" ;
		fco2_net_unc:_Endianness = "little" ;
	float fco2_para_unc(longitude, latitude, time) ;
		fco2_para_unc:units = "uatm" ;
		fco2_para_unc:long_name = "Fugacity of CO2 in seawater parameter uncertainty" ;
		fco2_para_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		fco2_para_unc:date_variable = "28/02/2025 17:28" ;
		fco2_para_unc:uncertainty_vals_lut = "[0.35, 0.4, 0.2, 0.1, 0.35, 0.4, 0.2, 0.1]" ;
		fco2_para_unc:uncertainty_vals_lut_parameters = "[\'CCI_SST_analysed_sst\', \'NOAA_ERSL_xCO2\', \'CCI_SSS_sss_CMEMS_so\', \'CMEMS_mlotst\', \'CCI_SST_analysed_sst_anom\', \'NOAA_ERSL_xCO2_anom\', \'CCI_SSS_sss_CMEMS_so_anom\', \'CMEMS_mlotst_anom\']" ;
		fco2_para_unc:lut_table_max_size = "20000" ;
		fco2_para_unc:_Storage = "contiguous" ;
		fco2_para_unc:_Endianness = "little" ;
	float latitude(latitude) ;
		latitude:units = "Degrees" ;
		latitude:standard_name = "Latitude" ;
		latitude:_Storage = "contiguous" ;
		latitude:_Endianness = "little" ;
	float longitude(longitude) ;
		longitude:units = "Degrees" ;
		longitude:standard_name = "Longitude" ;
		longitude:_Storage = "contiguous" ;
		longitude:_Endianness = "little" ;
	float time(time) ;
		time:units = "Days since 1970-01-15" ;
		time:standard_name = "Time of observations" ;
		time:_Storage = "contiguous" ;
		time:_Endianness = "little" ;
	float fco2_val_unc(longitude, latitude, time) ;
		fco2_val_unc:long_name = "Fugacity of CO2 in seawater evaluation uncertainty" ;
		fco2_val_unc:units = "uatm" ;
		fco2_val_unc:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		fco2_val_unc:date_generated = "28/02/2025 20:20" ;
		fco2_val_unc:_Storage = "contiguous" ;
		fco2_val_unc:_Endianness = "little" ;
	float fco2_tot_unc(longitude, latitude, time) ;
		fco2_tot_unc:date_generated = "28/02/2025 20:20" ;
		fco2_tot_unc:comment = "Combination offco2_val_unc, fco2_net_unc and fco2_para_unc in quadrature" ;
		fco2_tot_unc:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		fco2_tot_unc:units = "uatm" ;
		fco2_tot_unc:long_name = "Fugacity of CO2 in seawater total uncertainty" ;
		fco2_tot_unc:_Storage = "contiguous" ;
		fco2_tot_unc:_Endianness = "little" ;
	float flux(longitude, latitude, time) ;
		flux:units = "g C m-2 d-1" ;
		flux:calculations = "Flux calculations completed using FluxEngine" ;
		flux:long_name = "Air-sea CO2 flux" ;
		flux:comment = "Negative flux indicates atmosphere to ocean exchange" ;
		flux:date_generated = "01/03/2025 00:18" ;
		flux:_Storage = "contiguous" ;
		flux:_Endianness = "little" ;
	float flux_unc(longitude, latitude, time) ;
		flux_unc:long_name = "Air-sea CO2 flux total uncertainty" ;
		flux_unc:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc:seaice = "Sea ice uncertainty not included due to asymmetric nature of this flux uncertainty component" ;
		flux_unc:units = "Relative to flux" ;
		flux_unc:date_generated = "01/03/2025 00:18" ;
		flux_unc:_Storage = "contiguous" ;
		flux_unc:_Endianness = "little" ;
	float flux_unc_fco2sw(longitude, latitude, time) ;
		flux_unc_fco2sw:units = "Relative to flux" ;
		flux_unc_fco2sw:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_fco2sw:long_name = "Air-sea CO2 flux total fCO2sw uncertainty" ;
		flux_unc_fco2sw:date_generated = "01/03/2025 00:18" ;
		flux_unc_fco2sw:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_fco2sw:_Storage = "contiguous" ;
		flux_unc_fco2sw:_Endianness = "little" ;
	float flux_unc_fco2sw_net(longitude, latitude, time) ;
		flux_unc_fco2sw_net:units = "Relative to flux" ;
		flux_unc_fco2sw_net:date_generated = "01/03/2025 00:18" ;
		flux_unc_fco2sw_net:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_fco2sw_net:long_name = "Air-sea CO2 flux fCO2sw network uncertainty" ;
		flux_unc_fco2sw_net:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_fco2sw_net:_Storage = "contiguous" ;
		flux_unc_fco2sw_net:_Endianness = "little" ;
	float flux_unc_fco2sw_para(longitude, latitude, time) ;
		flux_unc_fco2sw_para:units = "Relative to flux" ;
		flux_unc_fco2sw_para:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_fco2sw_para:long_name = "Air-sea CO2 flux fCO2sw parameter uncertainty" ;
		flux_unc_fco2sw_para:date_generated = "01/03/2025 00:18" ;
		flux_unc_fco2sw_para:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_fco2sw_para:_Storage = "contiguous" ;
		flux_unc_fco2sw_para:_Endianness = "little" ;
	float flux_unc_fco2sw_val(longitude, latitude, time) ;
		flux_unc_fco2sw_val:units = "Relative to flux" ;
		flux_unc_fco2sw_val:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_fco2sw_val:long_name = "Air-sea CO2 flux fCO2sw evaluation uncertainty" ;
		flux_unc_fco2sw_val:date_generated = "01/03/2025 00:18" ;
		flux_unc_fco2sw_val:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_fco2sw_val:_Storage = "contiguous" ;
		flux_unc_fco2sw_val:_Endianness = "little" ;
	float flux_unc_k(longitude, latitude, time) ;
		flux_unc_k:long_name = "Air-sea CO2 flux gas transfer algorithm uncertainty" ;
		flux_unc_k:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_k:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_k:units = "Relative to flux" ;
		flux_unc_k:date_generated = "01/03/2025 00:18" ;
		flux_unc_k:fixed_value = "Algorithm uncertainty set at 20.0%" ;
		flux_unc_k:_Storage = "contiguous" ;
		flux_unc_k:_Endianness = "little" ;
	float flux_unc_wind(longitude, latitude, time) ;
		flux_unc_wind:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_wind:units = "Relative to flux" ;
		flux_unc_wind:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_wind:long_name = "Air-sea CO2 flux gas transfer uncertainty due to wind speed uncertainty" ;
		flux_unc_wind:date_generated = "01/03/2025 00:18" ;
		flux_unc_wind:_Storage = "contiguous" ;
		flux_unc_wind:_Endianness = "little" ;
	float flux_unc_schmidt(longitude, latitude, time) ;
		flux_unc_schmidt:units = "Relative to flux" ;
		flux_unc_schmidt:date_generated = "01/03/2025 00:18" ;
		flux_unc_schmidt:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_schmidt:long_name = "Air-sea CO2 flux Schmidt number uncertainty due to SST uncertainty" ;
		flux_unc_schmidt:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_schmidt:_Storage = "contiguous" ;
		flux_unc_schmidt:_Endianness = "little" ;
	float flux_unc_schmidt_fixed(longitude, latitude, time) ;
		flux_unc_schmidt_fixed:units = "Relative to flux" ;
		flux_unc_schmidt_fixed:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_schmidt_fixed:date_generated = "01/03/2025 00:18" ;
		flux_unc_schmidt_fixed:long_name = "Air-sea CO2 flux Schmidt number uncertainty due to algorithm uncertainty" ;
		flux_unc_schmidt_fixed:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_schmidt_fixed:_Storage = "contiguous" ;
		flux_unc_schmidt_fixed:_Endianness = "little" ;
	float flux_unc_ph2o(longitude, latitude, time) ;
		flux_unc_ph2o:units = "Relative to flux" ;
		flux_unc_ph2o:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_ph2o:long_name = "Air-sea CO2 flux pH2O correction uncertainty due to SST uncertainty" ;
		flux_unc_ph2o:date_generated = "01/03/2025 00:18" ;
		flux_unc_ph2o:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_ph2o:_Storage = "contiguous" ;
		flux_unc_ph2o:_Endianness = "little" ;
	float flux_unc_ph2o_fixed(longitude, latitude, time) ;
		flux_unc_ph2o_fixed:units = "Relative to flux" ;
		flux_unc_ph2o_fixed:date_generated = "01/03/2025 00:18" ;
		flux_unc_ph2o_fixed:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_ph2o_fixed:long_name = "Air-sea CO2 flux pH2O correction uncertainty due to algorithm uncertainty" ;
		flux_unc_ph2o_fixed:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_ph2o_fixed:_Storage = "contiguous" ;
		flux_unc_ph2o_fixed:_Endianness = "little" ;
	float flux_unc_xco2atm(longitude, latitude, time) ;
		flux_unc_xco2atm:units = "Relative to flux" ;
		flux_unc_xco2atm:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_xco2atm:long_name = "Air-sea CO2 flux xCO2atm uncertainty" ;
		flux_unc_xco2atm:date_generated = "01/03/2025 00:18" ;
		flux_unc_xco2atm:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_xco2atm:_Storage = "contiguous" ;
		flux_unc_xco2atm:_Endianness = "little" ;
	float flux_unc_solsubskin_unc(longitude, latitude, time) ;
		flux_unc_solsubskin_unc:units = "Relative to flux" ;
		flux_unc_solsubskin_unc:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_solsubskin_unc:long_name = "Air-sea CO2 flux subskin solubility uncertainty due to SST and SSS uncertainties" ;
		flux_unc_solsubskin_unc:date_generated = "01/03/2025 00:18" ;
		flux_unc_solsubskin_unc:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_solsubskin_unc:_Storage = "contiguous" ;
		flux_unc_solsubskin_unc:_Endianness = "little" ;
	float flux_unc_solsubskin_unc_fixed(longitude, latitude, time) ;
		flux_unc_solsubskin_unc_fixed:units = "Relative to flux" ;
		flux_unc_solsubskin_unc_fixed:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_solsubskin_unc_fixed:long_name = "Air-sea CO2 flux subskin solubility uncertainty due to algorithm uncertaintity" ;
		flux_unc_solsubskin_unc_fixed:date_generated = "01/03/2025 00:18" ;
		flux_unc_solsubskin_unc_fixed:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_solsubskin_unc_fixed:_Storage = "contiguous" ;
		flux_unc_solsubskin_unc_fixed:_Endianness = "little" ;
	float flux_unc_solskin_unc(longitude, latitude, time) ;
		flux_unc_solskin_unc:units = "Relative to flux" ;
		flux_unc_solskin_unc:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_solskin_unc:long_name = "Air-sea CO2 flux skin solubility uncertainty due to SST and SSS uncertainties" ;
		flux_unc_solskin_unc:date_generated = "01/03/2025 00:18" ;
		flux_unc_solskin_unc:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_solskin_unc:_Storage = "contiguous" ;
		flux_unc_solskin_unc:_Endianness = "little" ;
	float flux_unc_solskin_unc_fixed(longitude, latitude, time) ;
		flux_unc_solskin_unc_fixed:units = "Relative to flux" ;
		flux_unc_solskin_unc_fixed:comment = "Multiple by absolute flux to get uncertainty in g C m-2 d-1" ;
		flux_unc_solskin_unc_fixed:long_name = "Air-sea CO2 flux skin solubility uncertainty due to algorithm uncertaintity" ;
		flux_unc_solskin_unc_fixed:date_generated = "01/03/2025 00:18" ;
		flux_unc_solskin_unc_fixed:uncertainties = "Uncertainties considered 95% confidence (2 sigma)" ;
		flux_unc_solskin_unc_fixed:_Storage = "contiguous" ;
		flux_unc_solskin_unc_fixed:_Endianness = "little" ;
	float ice(longitude, latitude, time) ;
		ice:units = "Proportion" ;
		ice:long_name = "Proportion of ice cover" ;
		ice:comment = "See the OceanICU framework config file for the ice dataset used in these calculations" ;
		ice:date_generated = "01/03/2025 00:18" ;
		ice:_Storage = "contiguous" ;
		ice:_Endianness = "little" ;
	float subskin_temp(longitude, latitude, time) ;
		subskin_temp:units = "Kelvin" ;
		subskin_temp:long_name = "Subskin temperature" ;
		subskin_temp:date_generated = "01/03/2025 00:18" ;
		subskin_temp:comment = "See the OceanICU framework config file for the SST subskin dataset used in these calculations" ;
		subskin_temp:_Storage = "contiguous" ;
		subskin_temp:_Endianness = "little" ;
	float skin_temp(longitude, latitude, time) ;
		skin_temp:units = "Kelvin" ;
		skin_temp:long_name = "Skin temperature" ;
		skin_temp:comment = "See the OceanICU framework config file for the SST skin dataset used in these calculations" ;
		skin_temp:date_generated = "01/03/2025 00:18" ;
		skin_temp:_Storage = "contiguous" ;
		skin_temp:_Endianness = "little" ;
	float skin_salinity(longitude, latitude, time) ;
		skin_salinity:units = "psu" ;
		skin_salinity:long_name = "Skin salinity" ;
		skin_salinity:comment = "See the OceanICU framework config file for the SSS skin dataset used in these calculations" ;
		skin_salinity:date_generated = "01/03/2025 00:18" ;
		skin_salinity:_Storage = "contiguous" ;
		skin_salinity:_Endianness = "little" ;
	float subskin_salinity(longitude, latitude, time) ;
		subskin_salinity:units = "psu" ;
		subskin_salinity:long_name = "Subskin salinity" ;
		subskin_salinity:comment = "See the OceanICU framework config file for the SSS subskin dataset used in these calculations" ;
		subskin_salinity:date_generated = "01/03/2025 00:18" ;
		subskin_salinity:_Storage = "contiguous" ;
		subskin_salinity:_Endianness = "little" ;
	float ta(longitude, latitude, time) ;
		ta:units = "umol/kg" ;
		ta:long_name = "Total Alkalinity" ;
		ta:comment = "" ;
		ta:date_variable = "02/03/2025 11:27" ;
		ta:_Storage = "contiguous" ;
		ta:_Endianness = "little" ;
	float ta_net_unc(longitude, latitude, time) ;
		ta_net_unc:units = "umol/kg" ;
		ta_net_unc:long_name = "Total Alkalinity network uncertainty" ;
		ta_net_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		ta_net_unc:date_variable = "02/03/2025 11:27" ;
		ta_net_unc:_Storage = "contiguous" ;
		ta_net_unc:_Endianness = "little" ;
	float ta_tot_unc(longitude, latitude, time) ;
		ta_tot_unc:units = "umol/kg" ;
		ta_tot_unc:long_name = "Total Alkalinity total uncertainty" ;
		ta_tot_unc:comment = "Combination ofta_val_unc, ta_net_unc and ta_para_unc in quadrature" ;
		ta_tot_unc:date_variable = "02/03/2025 11:27" ;
		ta_tot_unc:_Storage = "contiguous" ;
		ta_tot_unc:_Endianness = "little" ;
	float ta_val_unc(longitude, latitude, time) ;
		ta_val_unc:comment = "" ;
		ta_val_unc:units = "umol/kg" ;
		ta_val_unc:long_name = "Total Alkalinity evaluation uncertainty" ;
		ta_val_unc:date_variable = "02/03/2025 11:27" ;
		ta_val_unc:_Storage = "contiguous" ;
		ta_val_unc:_Endianness = "little" ;
	float ta_para_unc(longitude, latitude, time) ;
		ta_para_unc:units = "umol/kg" ;
		ta_para_unc:long_name = "Total Alkalinity parameter uncertainty" ;
		ta_para_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		ta_para_unc:date_variable = "02/03/2025 11:27" ;
		ta_para_unc:_Storage = "contiguous" ;
		ta_para_unc:_Endianness = "little" ;
	float dic(longitude, latitude, time) ;
		dic:units = "umol/kg" ;
		dic:long_name = "Dissolved Inorganic Carbon in seawater" ;
		dic:comment = "" ;
		dic:date_variable = "02/03/2025 13:59" ;
		dic:_Storage = "contiguous" ;
		dic:_Endianness = "little" ;
	float dic_tot_unc(longitude, latitude, time) ;
		dic_tot_unc:units = "umol/kg" ;
		dic_tot_unc:long_name = "Dissolved Inorganic Carbon in seawater total uncertainty" ;
		dic_tot_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		dic_tot_unc:date_variable = "02/03/2025 13:59" ;
		dic_tot_unc:_Storage = "contiguous" ;
		dic_tot_unc:_Endianness = "little" ;
	float dic_ta_unc(longitude, latitude, time) ;
		dic_ta_unc:units = "umol/kg" ;
		dic_ta_unc:long_name = "Dissolved Inorganic Carbon in seawater alkalinity uncertainty" ;
		dic_ta_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		dic_ta_unc:date_variable = "02/03/2025 13:59" ;
		dic_ta_unc:_Storage = "contiguous" ;
		dic_ta_unc:_Endianness = "little" ;
	float dic_fco2_unc(longitude, latitude, time) ;
		dic_fco2_unc:units = "umol/kg" ;
		dic_fco2_unc:long_name = "Dissolved Inorganic Carbon in seawater fCO2(sw) uncertainty" ;
		dic_fco2_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		dic_fco2_unc:date_variable = "02/03/2025 13:59" ;
		dic_fco2_unc:_Storage = "contiguous" ;
		dic_fco2_unc:_Endianness = "little" ;
	float dic_sst_unc(longitude, latitude, time) ;
		dic_sst_unc:units = "umol/kg" ;
		dic_sst_unc:long_name = "Dissolved Inorganic Carbon in seawater SST uncertainty" ;
		dic_sst_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		dic_sst_unc:date_variable = "02/03/2025 13:59" ;
		dic_sst_unc:_Storage = "contiguous" ;
		dic_sst_unc:_Endianness = "little" ;
	float dic_sss_unc(longitude, latitude, time) ;
		dic_sss_unc:units = "umol/kg" ;
		dic_sss_unc:long_name = "Dissolved Inorganic Carbon in seawater SSS uncertainty" ;
		dic_sss_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		dic_sss_unc:date_variable = "02/03/2025 13:59" ;
		dic_sss_unc:_Storage = "contiguous" ;
		dic_sss_unc:_Endianness = "little" ;
	float dic_phos_unc(longitude, latitude, time) ;
		dic_phos_unc:units = "umol/kg" ;
		dic_phos_unc:date_variable = "02/03/2025 13:59" ;
		dic_phos_unc:long_name = "Dissolved Inorganic Carbon in seawater phosphate uncertainty" ;
		dic_phos_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		dic_phos_unc:_Storage = "contiguous" ;
		dic_phos_unc:_Endianness = "little" ;
	float dic_sili_unc(longitude, latitude, time) ;
		dic_sili_unc:units = "umol/kg" ;
		dic_sili_unc:long_name = "Dissolved Inorganic Carbon in seawater silicate uncertainty" ;
		dic_sili_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		dic_sili_unc:date_variable = "02/03/2025 13:59" ;
		dic_sili_unc:_Storage = "contiguous" ;
		dic_sili_unc:_Endianness = "little" ;
	float pH(longitude, latitude, time) ;
		pH:comment = "" ;
		pH:units = "-log([H+])" ;
		pH:long_name = "pH on total scale" ;
		pH:date_variable = "02/03/2025 13:59" ;
		pH:_Storage = "contiguous" ;
		pH:_Endianness = "little" ;
	float pH_tot_unc(longitude, latitude, time) ;
		pH_tot_unc:units = "-log([H+])" ;
		pH_tot_unc:date_variable = "02/03/2025 13:59" ;
		pH_tot_unc:long_name = "pH on total scale total uncertainty" ;
		pH_tot_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		pH_tot_unc:_Storage = "contiguous" ;
		pH_tot_unc:_Endianness = "little" ;
	float pH_ta_unc(longitude, latitude, time) ;
		pH_ta_unc:units = "-log([H+])" ;
		pH_ta_unc:date_variable = "02/03/2025 13:59" ;
		pH_ta_unc:long_name = "pH on total scale alkalinity uncertainty" ;
		pH_ta_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		pH_ta_unc:_Storage = "contiguous" ;
		pH_ta_unc:_Endianness = "little" ;
	float pH_fco2_unc(longitude, latitude, time) ;
		pH_fco2_unc:units = "-log([H+])" ;
		pH_fco2_unc:long_name = "pH on total scale fCO2(sw) uncertainty" ;
		pH_fco2_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		pH_fco2_unc:date_variable = "02/03/2025 13:59" ;
		pH_fco2_unc:_Storage = "contiguous" ;
		pH_fco2_unc:_Endianness = "little" ;
	float pH_sst_unc(longitude, latitude, time) ;
		pH_sst_unc:units = "-log([H+])" ;
		pH_sst_unc:long_name = "pH on total scale SST uncertainty" ;
		pH_sst_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		pH_sst_unc:date_variable = "02/03/2025 13:59" ;
		pH_sst_unc:_Storage = "contiguous" ;
		pH_sst_unc:_Endianness = "little" ;
	float pH_sss_unc(longitude, latitude, time) ;
		pH_sss_unc:units = "-log([H+])" ;
		pH_sss_unc:long_name = "pH on total scale SSS uncertainty" ;
		pH_sss_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		pH_sss_unc:date_variable = "02/03/2025 13:59" ;
		pH_sss_unc:_Storage = "contiguous" ;
		pH_sss_unc:_Endianness = "little" ;
	float pH_phos_unc(longitude, latitude, time) ;
		pH_phos_unc:units = "-log([H+])" ;
		pH_phos_unc:long_name = "pH on total scale phosphate uncertainty" ;
		pH_phos_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		pH_phos_unc:date_variable = "02/03/2025 13:59" ;
		pH_phos_unc:_Storage = "contiguous" ;
		pH_phos_unc:_Endianness = "little" ;
	float pH_sili_unc(longitude, latitude, time) ;
		pH_sili_unc:units = "-log([H+])" ;
		pH_sili_unc:long_name = "pH on total scale silicate uncertainty" ;
		pH_sili_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		pH_sili_unc:date_variable = "02/03/2025 13:59" ;
		pH_sili_unc:_Storage = "contiguous" ;
		pH_sili_unc:_Endianness = "little" ;
	float saturation_aragonite(longitude, latitude, time) ;
		saturation_aragonite:units = "unitless" ;
		saturation_aragonite:long_name = "Saturation state of Aragonite" ;
		saturation_aragonite:comment = "" ;
		saturation_aragonite:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite:_Storage = "contiguous" ;
		saturation_aragonite:_Endianness = "little" ;
	float saturation_aragonite_tot_unc(longitude, latitude, time) ;
		saturation_aragonite_tot_unc:units = "unitless" ;
		saturation_aragonite_tot_unc:long_name = "Saturation state of Aragonite total uncertainty" ;
		saturation_aragonite_tot_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		saturation_aragonite_tot_unc:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite_tot_unc:_Storage = "contiguous" ;
		saturation_aragonite_tot_unc:_Endianness = "little" ;
	float saturation_aragonite_ta_unc(longitude, latitude, time) ;
		saturation_aragonite_ta_unc:units = "unitless" ;
		saturation_aragonite_ta_unc:long_name = "Saturation state of Aragonite alkalinity uncertainty" ;
		saturation_aragonite_ta_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		saturation_aragonite_ta_unc:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite_ta_unc:_Storage = "contiguous" ;
		saturation_aragonite_ta_unc:_Endianness = "little" ;
	float saturation_aragonite_fco2_unc(longitude, latitude, time) ;
		saturation_aragonite_fco2_unc:units = "unitless" ;
		saturation_aragonite_fco2_unc:long_name = "Saturation state of Aragonite fCO2(sw) uncertainty" ;
		saturation_aragonite_fco2_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		saturation_aragonite_fco2_unc:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite_fco2_unc:_Storage = "contiguous" ;
		saturation_aragonite_fco2_unc:_Endianness = "little" ;
	float saturation_aragonite_sst_unc(longitude, latitude, time) ;
		saturation_aragonite_sst_unc:units = "unitless" ;
		saturation_aragonite_sst_unc:long_name = "Saturation state of Aragonite SST uncertainty" ;
		saturation_aragonite_sst_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		saturation_aragonite_sst_unc:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite_sst_unc:_Storage = "contiguous" ;
		saturation_aragonite_sst_unc:_Endianness = "little" ;
	float saturation_aragonite_sss_unc(longitude, latitude, time) ;
		saturation_aragonite_sss_unc:units = "unitless" ;
		saturation_aragonite_sss_unc:long_name = "Saturation state of Aragonite SSS uncertainty" ;
		saturation_aragonite_sss_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		saturation_aragonite_sss_unc:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite_sss_unc:_Storage = "contiguous" ;
		saturation_aragonite_sss_unc:_Endianness = "little" ;
	float saturation_aragonite_phos_unc(longitude, latitude, time) ;
		saturation_aragonite_phos_unc:units = "unitless" ;
		saturation_aragonite_phos_unc:long_name = "Saturation state of Aragonite phosphate uncertainty" ;
		saturation_aragonite_phos_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		saturation_aragonite_phos_unc:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite_phos_unc:_Storage = "contiguous" ;
		saturation_aragonite_phos_unc:_Endianness = "little" ;
	float saturation_aragonite_sili_unc(longitude, latitude, time) ;
		saturation_aragonite_sili_unc:units = "unitless" ;
		saturation_aragonite_sili_unc:long_name = "Saturation state of Aragonite silicate uncertainty" ;
		saturation_aragonite_sili_unc:comment = "Uncertainties considered 95% confidence (2 sigma)" ;
		saturation_aragonite_sili_unc:date_variable = "02/03/2025 13:59" ;
		saturation_aragonite_sili_unc:_Storage = "contiguous" ;
		saturation_aragonite_sili_unc:_Endianness = "little" ;

// global attributes:
		:date_file_generated = "28/02/2025 17:28" ;
		:code_by = "Daniel J. Ford (d.ford@exeter.ac.uk)" ;
		:code_location = "https://github.com/JamieLab/OceanICU" ;
		:_NCProperties = "version=2,netcdf=4.9.2,hdf5=1.14.4" ;
		:_SuperblockVersion = 2 ;
		:_IsNetcdf4 = 0 ;
		:_Format = "netCDF-4 classic model" ;
}
