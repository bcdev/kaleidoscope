netcdf mercatorglorys12v1_gl12_mean_200001 {
dimensions:
	longitude = 4320 ;
	latitude = 2041 ;
	depth = 50 ;
	time = 1 ;
variables:
	float longitude(longitude) ;
		longitude:_FillValue = NaNf ;
		longitude:valid_min = -180.f ;
		longitude:valid_max = 179.9167f ;
		longitude:step = 0.08332825f ;
		longitude:units = "degrees_east" ;
		longitude:unit_long = "Degrees East" ;
		longitude:long_name = "Longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:axis = "X" ;
		longitude:_Storage = "chunked" ;
		longitude:_ChunkSizes = 4320 ;
		longitude:_DeflateLevel = 1 ;
		longitude:_Endianness = "little" ;
	float latitude(latitude) ;
		latitude:_FillValue = NaNf ;
		latitude:valid_min = -80.f ;
		latitude:valid_max = 90.f ;
		latitude:step = 0.08333588f ;
		latitude:units = "degrees_north" ;
		latitude:unit_long = "Degrees North" ;
		latitude:long_name = "Latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:axis = "Y" ;
		latitude:_Storage = "chunked" ;
		latitude:_ChunkSizes = 2041 ;
		latitude:_DeflateLevel = 1 ;
		latitude:_Endianness = "little" ;
	float depth(depth) ;
		depth:_FillValue = NaNf ;
		depth:valid_min = 0.494025f ;
		depth:valid_max = 5727.917f ;
		depth:units = "m" ;
		depth:positive = "down" ;
		depth:unit_long = "Meters" ;
		depth:long_name = "Depth" ;
		depth:standard_name = "depth" ;
		depth:axis = "Z" ;
		depth:_Storage = "chunked" ;
		depth:_ChunkSizes = 50 ;
		depth:_DeflateLevel = 1 ;
		depth:_Endianness = "little" ;
	short mlotst(time, latitude, longitude) ;
		mlotst:_FillValue = -32767s ;
		mlotst:long_name = "Density ocean mixed layer thickness" ;
		mlotst:standard_name = "ocean_mixed_layer_thickness_defined_by_sigma_theta" ;
		mlotst:units = "m" ;
		mlotst:unit_long = "Meters" ;
		mlotst:valid_min = 1s ;
		mlotst:valid_max = 8881s ;
		mlotst:cell_methods = "area: mean" ;
		mlotst:add_offset = -0.152592554688454 ;
		mlotst:scale_factor = 0.152592554688454 ;
		mlotst:_Storage = "chunked" ;
		mlotst:_ChunkSizes = 1, 1021, 2160 ;
		mlotst:_DeflateLevel = 1 ;
		mlotst:_Endianness = "little" ;
	short zos(time, latitude, longitude) ;
		zos:_FillValue = -32767s ;
		zos:long_name = "Sea surface height" ;
		zos:standard_name = "sea_surface_height_above_geoid" ;
		zos:units = "m" ;
		zos:unit_long = "Meters" ;
		zos:valid_min = -6382s ;
		zos:valid_max = 4883s ;
		zos:cell_methods = "area: mean" ;
		zos:add_offset = 0. ;
		zos:scale_factor = 0.000305185094475746 ;
		zos:_Storage = "chunked" ;
		zos:_ChunkSizes = 1, 1021, 2160 ;
		zos:_DeflateLevel = 1 ;
		zos:_Endianness = "little" ;
	short bottomT(time, latitude, longitude) ;
		bottomT:_FillValue = -32767s ;
		bottomT:long_name = "Sea floor potential temperature" ;
		bottomT:standard_name = "sea_water_potential_temperature_at_sea_floor" ;
		bottomT:units = "degrees_C" ;
		bottomT:unit_long = "Degrees Celsius" ;
		bottomT:valid_min = -32639s ;
		bottomT:valid_max = 18498s ;
		bottomT:cell_methods = "area: mean" ;
		bottomT:add_offset = 21. ;
		bottomT:scale_factor = 0.000732444226741791 ;
		bottomT:_Storage = "chunked" ;
		bottomT:_ChunkSizes = 1, 1021, 2160 ;
		bottomT:_DeflateLevel = 1 ;
		bottomT:_Endianness = "little" ;
	short sithick(time, latitude, longitude) ;
		sithick:_FillValue = -32767s ;
		sithick:long_name = "Sea ice thickness" ;
		sithick:standard_name = "sea_ice_thickness" ;
		sithick:units = "m" ;
		sithick:unit_long = "Meters" ;
		sithick:valid_min = 1s ;
		sithick:valid_max = 8041s ;
		sithick:cell_methods = "area: mean where sea_ice" ;
		sithick:add_offset = -0.000762962736189365 ;
		sithick:scale_factor = 0.000762962736189365 ;
		sithick:_Storage = "chunked" ;
		sithick:_ChunkSizes = 1, 1021, 2160 ;
		sithick:_DeflateLevel = 1 ;
		sithick:_Endianness = "little" ;
	short siconc(time, latitude, longitude) ;
		siconc:_FillValue = -32767s ;
		siconc:long_name = "Ice concentration" ;
		siconc:standard_name = "sea_ice_area_fraction" ;
		siconc:units = "1" ;
		siconc:unit_long = "Fraction" ;
		siconc:valid_min = 1s ;
		siconc:valid_max = 28317s ;
		siconc:cell_methods = "area: mean where sea_ice" ;
		siconc:add_offset = -3.81481368094683e-05 ;
		siconc:scale_factor = 3.81481368094683e-05 ;
		siconc:_Storage = "chunked" ;
		siconc:_ChunkSizes = 1, 1021, 2160 ;
		siconc:_DeflateLevel = 1 ;
		siconc:_Endianness = "little" ;
	short usi(time, latitude, longitude) ;
		usi:_FillValue = -32767s ;
		usi:long_name = "Sea ice eastward velocity" ;
		usi:standard_name = "eastward_sea_ice_velocity" ;
		usi:units = "m s-1" ;
		usi:unit_long = "Meters per second" ;
		usi:valid_min = -20539s ;
		usi:valid_max = 32652s ;
		usi:cell_methods = "area: mean where sea_ice" ;
		usi:add_offset = 0. ;
		usi:scale_factor = 3.05185094475746e-05 ;
		usi:_Storage = "chunked" ;
		usi:_ChunkSizes = 1, 1021, 2160 ;
		usi:_DeflateLevel = 1 ;
		usi:_Endianness = "little" ;
	short vsi(time, latitude, longitude) ;
		vsi:_FillValue = -32767s ;
		vsi:long_name = "Sea ice northward velocity" ;
		vsi:standard_name = "northward_sea_ice_velocity" ;
		vsi:units = "m s-1" ;
		vsi:unit_long = "Meters per second" ;
		vsi:valid_min = -32637s ;
		vsi:valid_max = 24967s ;
		vsi:cell_methods = "area: mean where sea_ice" ;
		vsi:add_offset = 0. ;
		vsi:scale_factor = 3.05185094475746e-05 ;
		vsi:_Storage = "chunked" ;
		vsi:_ChunkSizes = 1, 1021, 2160 ;
		vsi:_DeflateLevel = 1 ;
		vsi:_Endianness = "little" ;
	short thetao(time, depth, latitude, longitude) ;
		thetao:_FillValue = -32767s ;
		thetao:long_name = "Temperature" ;
		thetao:standard_name = "sea_water_potential_temperature" ;
		thetao:units = "degrees_C" ;
		thetao:unit_long = "Degrees Celsius" ;
		thetao:valid_min = -32764s ;
		thetao:valid_max = 18468s ;
		thetao:cell_methods = "area: mean" ;
		thetao:add_offset = 21. ;
		thetao:scale_factor = 0.000732444226741791 ;
		thetao:_Storage = "chunked" ;
		thetao:_ChunkSizes = 1, 10, 511, 1080 ;
		thetao:_DeflateLevel = 1 ;
		thetao:_Endianness = "little" ;
	short so(time, depth, latitude, longitude) ;
		so:_FillValue = -32767s ;
		so:long_name = "Salinity" ;
		so:standard_name = "sea_water_salinity" ;
		so:units = "1e-3" ;
		so:unit_long = "Practical Salinity Unit" ;
		so:valid_min = 1s ;
		so:valid_max = 27353s ;
		so:cell_methods = "area: mean" ;
		so:add_offset = -0.00152592547237873 ;
		so:scale_factor = 0.00152592547237873 ;
		so:_Storage = "chunked" ;
		so:_ChunkSizes = 1, 10, 511, 1080 ;
		so:_DeflateLevel = 1 ;
		so:_Endianness = "little" ;
	short uo(time, depth, latitude, longitude) ;
		uo:_FillValue = -32767s ;
		uo:long_name = "Eastward velocity" ;
		uo:standard_name = "eastward_sea_water_velocity" ;
		uo:units = "m s-1" ;
		uo:unit_long = "Meters per second" ;
		uo:valid_min = -3510s ;
		uo:valid_max = 3894s ;
		uo:cell_methods = "area: mean" ;
		uo:add_offset = 0. ;
		uo:scale_factor = 0.000610370188951492 ;
		uo:_Storage = "chunked" ;
		uo:_ChunkSizes = 1, 10, 511, 1080 ;
		uo:_DeflateLevel = 1 ;
		uo:_Endianness = "little" ;
	short vo(time, depth, latitude, longitude) ;
		vo:_FillValue = -32767s ;
		vo:long_name = "Northward velocity" ;
		vo:standard_name = "northward_sea_water_velocity" ;
		vo:units = "m s-1" ;
		vo:unit_long = "Meters per second" ;
		vo:valid_min = -3234s ;
		vo:valid_max = 3332s ;
		vo:cell_methods = "area: mean" ;
		vo:add_offset = 0. ;
		vo:scale_factor = 0.000610370188951492 ;
		vo:_Storage = "chunked" ;
		vo:_ChunkSizes = 1, 10, 511, 1080 ;
		vo:_DeflateLevel = 1 ;
		vo:_Endianness = "little" ;
	double time(time) ;
		time:_FillValue = NaN ;
		time:units = "hours since 1950-01-01" ;
		time:axis = "T" ;
		time:long_name = "Time (hours since 1950-01-01)" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
		time:_Storage = "chunked" ;
		time:_ChunkSizes = 1 ;
		time:_DeflateLevel = 1 ;
		time:_Endianness = "little" ;

// global attributes:
		:title = "Monthly mean fields for product GLOBAL_REANALYSIS_PHY_001_030" ;
		:references = "http://marine.copernicus.eu" ;
		:credit = "E.U. Copernicus Marine Service Information (CMEMS)" ;
		:licence = "http://marine.copernicus.eu/services-portfolio/service-commitments-and-licence/" ;
		:contact = "servicedesk.cmems@mercator-ocean.eu" ;
		:producer = "CMEMS - Global Monitoring and Forecasting Centre" ;
		:institution = "Mercator Ocean" ;
		:Conventions = "CF-1.6" ;
		:area = "GLOBAL" ;
		:product = "GLOBAL_REANALYSIS_001_030" ;
		:dataset = "global-reanalysis-001-030-monthly" ;
		:source = "MERCATOR GLORYS12V1" ;
		:product_user_manual = "http://marine.copernicus.eu/documents/PUM/CMEMS-GLO-PUM-001-030.pdf" ;
		:quality_information_document = "http://marine.copernicus.eu/documents/QUID/CMEMS-GLO-QUID-001-030.pdf" ;
		:_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.18" ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
}
